module picorv32a (clk,
    mem_instr,
    mem_la_read,
    mem_la_write,
    mem_ready,
    mem_valid,
    pcpi_ready,
    pcpi_valid,
    pcpi_wait,
    pcpi_wr,
    resetn,
    trace_valid,
    trap,
    VPWR,
    VGND,
    eoi,
    irq,
    mem_addr,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    mem_rdata,
    mem_wdata,
    mem_wstrb,
    pcpi_insn,
    pcpi_rd,
    pcpi_rs1,
    pcpi_rs2,
    trace_data);
 input clk;
 output mem_instr;
 output mem_la_read;
 output mem_la_write;
 input mem_ready;
 output mem_valid;
 input pcpi_ready;
 output pcpi_valid;
 input pcpi_wait;
 input pcpi_wr;
 input resetn;
 output trace_valid;
 output trap;
 input VPWR;
 input VGND;
 output [31:0] eoi;
 input [31:0] irq;
 output [31:0] mem_addr;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 output [31:0] pcpi_insn;
 input [31:0] pcpi_rd;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 output [35:0] trace_data;

 sky130_fd_sc_hd__and2_2 _15294_ (.A(net237),
    .B(net65),
    .X(_12629_));
 sky130_fd_sc_hd__and2_1 _15295_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .X(_12630_));
 sky130_fd_sc_hd__buf_2 _15296_ (.A(\mem_state[0] ),
    .X(_12631_));
 sky130_fd_sc_hd__nor2_8 _15297_ (.A(\mem_state[1] ),
    .B(_12631_),
    .Y(_00290_));
 sky130_fd_sc_hd__o21ba_4 _15298_ (.A1(_12629_),
    .A2(_12630_),
    .B1_N(_00290_),
    .X(_12632_));
 sky130_vsdinv _15299_ (.A(net237),
    .Y(_12633_));
 sky130_vsdinv _15300_ (.A(net65),
    .Y(_12634_));
 sky130_fd_sc_hd__nor2_8 _15301_ (.A(mem_do_wdata),
    .B(mem_do_rdata),
    .Y(_12635_));
 sky130_vsdinv _15302_ (.A(mem_do_rinst),
    .Y(_12636_));
 sky130_fd_sc_hd__o31ai_1 _15303_ (.A1(_12633_),
    .A2(_12634_),
    .A3(_12635_),
    .B1(_12636_),
    .Y(_12637_));
 sky130_fd_sc_hd__clkbuf_4 _15304_ (.A(net101),
    .X(_12638_));
 sky130_fd_sc_hd__nand3_4 _15305_ (.A(_12632_),
    .B(net456),
    .C(_12638_),
    .Y(_12639_));
 sky130_fd_sc_hd__clkbuf_4 _15306_ (.A(mem_do_prefetch),
    .X(_12640_));
 sky130_vsdinv _15307_ (.A(net101),
    .Y(_12641_));
 sky130_fd_sc_hd__buf_2 _15308_ (.A(_12641_),
    .X(_12642_));
 sky130_fd_sc_hd__buf_4 _15309_ (.A(_12642_),
    .X(_12643_));
 sky130_fd_sc_hd__a21oi_4 _15310_ (.A1(_12639_),
    .A2(_12640_),
    .B1(_12643_),
    .Y(_12644_));
 sky130_fd_sc_hd__clkbuf_2 _15311_ (.A(mem_do_rdata),
    .X(_12645_));
 sky130_fd_sc_hd__and2_1 _15312_ (.A(_12645_),
    .B(\cpu_state[6] ),
    .X(_12646_));
 sky130_fd_sc_hd__clkbuf_2 _15313_ (.A(_12646_),
    .X(_00319_));
 sky130_fd_sc_hd__a21oi_2 _15314_ (.A1(_12644_),
    .A2(_00319_),
    .B1(_00332_),
    .Y(_12647_));
 sky130_fd_sc_hd__clkbuf_2 _15315_ (.A(_12638_),
    .X(_12648_));
 sky130_fd_sc_hd__clkbuf_4 _15316_ (.A(_12648_),
    .X(_12649_));
 sky130_fd_sc_hd__buf_4 _15317_ (.A(_12649_),
    .X(_12650_));
 sky130_fd_sc_hd__clkbuf_2 _15318_ (.A(\cpu_state[6] ),
    .X(_12651_));
 sky130_fd_sc_hd__buf_2 _15319_ (.A(_12651_),
    .X(_12652_));
 sky130_fd_sc_hd__a221o_1 _15320_ (.A1(instr_lb),
    .A2(_12652_),
    .B1(_12644_),
    .B2(_00319_),
    .C1(_00332_),
    .X(_12653_));
 sky130_fd_sc_hd__o211a_1 _15321_ (.A1(latched_is_lb),
    .A2(_12647_),
    .B1(_12650_),
    .C1(_12653_),
    .X(_04071_));
 sky130_fd_sc_hd__buf_4 _15322_ (.A(_12648_),
    .X(_12654_));
 sky130_fd_sc_hd__buf_1 _15323_ (.A(_12654_),
    .X(_12655_));
 sky130_fd_sc_hd__buf_4 _15324_ (.A(_12655_),
    .X(_12656_));
 sky130_vsdinv _15325_ (.A(instr_lh),
    .Y(_12657_));
 sky130_vsdinv _15326_ (.A(\cpu_state[6] ),
    .Y(_12658_));
 sky130_fd_sc_hd__buf_2 _15327_ (.A(_12658_),
    .X(_12659_));
 sky130_fd_sc_hd__buf_4 _15328_ (.A(_12659_),
    .X(_12660_));
 sky130_fd_sc_hd__o21ai_1 _15329_ (.A1(_12657_),
    .A2(_12660_),
    .B1(_12647_),
    .Y(_12661_));
 sky130_fd_sc_hd__o211a_1 _15330_ (.A1(latched_is_lh),
    .A2(_12647_),
    .B1(_12656_),
    .C1(_12661_),
    .X(_04070_));
 sky130_fd_sc_hd__and2b_1 _15331_ (.A_N(instr_retirq),
    .B(\cpu_state[2] ),
    .X(_12662_));
 sky130_fd_sc_hd__clkbuf_4 _15332_ (.A(latched_branch),
    .X(_12663_));
 sky130_fd_sc_hd__o21bai_1 _15333_ (.A1(_00331_),
    .A2(_12662_),
    .B1_N(_12663_),
    .Y(_12664_));
 sky130_fd_sc_hd__o311a_1 _15334_ (.A1(_15243_),
    .A2(_00331_),
    .A3(_12662_),
    .B1(_12650_),
    .C1(_12664_),
    .X(_04069_));
 sky130_vsdinv _15335_ (.A(\mem_state[1] ),
    .Y(_12665_));
 sky130_fd_sc_hd__buf_4 _15336_ (.A(mem_do_rinst),
    .X(_12666_));
 sky130_fd_sc_hd__and2_1 _15337_ (.A(_12631_),
    .B(_12666_),
    .X(_12667_));
 sky130_fd_sc_hd__and3b_1 _15338_ (.A_N(_12631_),
    .B(net237),
    .C(net65),
    .X(_12668_));
 sky130_vsdinv _15339_ (.A(net408),
    .Y(_12669_));
 sky130_fd_sc_hd__nor2_8 _15340_ (.A(_12666_),
    .B(mem_do_prefetch),
    .Y(_12670_));
 sky130_fd_sc_hd__nand3_2 _15341_ (.A(_00290_),
    .B(_12635_),
    .C(_12670_),
    .Y(_12671_));
 sky130_fd_sc_hd__o311ai_4 _15342_ (.A1(_12665_),
    .A2(_12667_),
    .A3(_12668_),
    .B1(_12669_),
    .C1(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__a21boi_4 _15343_ (.A1(_12672_),
    .A2(_12649_),
    .B1_N(_00300_),
    .Y(_12673_));
 sky130_fd_sc_hd__clkbuf_4 _15344_ (.A(_12638_),
    .X(_12674_));
 sky130_fd_sc_hd__nor2b_4 _15345_ (.A(net408),
    .B_N(_12674_),
    .Y(_12675_));
 sky130_fd_sc_hd__clkbuf_2 _15346_ (.A(_12675_),
    .X(_12676_));
 sky130_fd_sc_hd__nand3_1 _15347_ (.A(_12673_),
    .B(_15208_),
    .C(_12676_),
    .Y(_12677_));
 sky130_fd_sc_hd__o21ai_1 _15348_ (.A1(_12665_),
    .A2(_12673_),
    .B1(_12677_),
    .Y(_04068_));
 sky130_vsdinv _15349_ (.A(_12631_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand3_1 _15350_ (.A(_12673_),
    .B(_15207_),
    .C(_12676_),
    .Y(_12679_));
 sky130_fd_sc_hd__o21ai_1 _15351_ (.A1(_12678_),
    .A2(_12673_),
    .B1(_12679_),
    .Y(_04067_));
 sky130_fd_sc_hd__nor2_4 _15352_ (.A(_12636_),
    .B(_12639_),
    .Y(_12680_));
 sky130_fd_sc_hd__buf_2 _15353_ (.A(_12680_),
    .X(_12681_));
 sky130_fd_sc_hd__clkbuf_4 _15354_ (.A(_12681_),
    .X(_15210_));
 sky130_fd_sc_hd__inv_2 _15355_ (.A(\decoded_rs1[4] ),
    .Y(_00366_));
 sky130_vsdinv _15356_ (.A(_00327_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand3b_4 _15357_ (.A_N(_00326_),
    .B(_00325_),
    .C(_00324_),
    .Y(_12683_));
 sky130_vsdinv _15358_ (.A(_00329_),
    .Y(_12684_));
 sky130_vsdinv _15359_ (.A(_00328_),
    .Y(_12685_));
 sky130_vsdinv _15360_ (.A(_00330_),
    .Y(_12686_));
 sky130_fd_sc_hd__nand3_1 _15361_ (.A(_12684_),
    .B(_12685_),
    .C(_12686_),
    .Y(_12687_));
 sky130_fd_sc_hd__or4_4 _15362_ (.A(\mem_rdata_latched[28] ),
    .B(_12682_),
    .C(_12683_),
    .D(_12687_),
    .X(_12688_));
 sky130_fd_sc_hd__or3_1 _15363_ (.A(\mem_rdata_latched[31] ),
    .B(\mem_rdata_latched[30] ),
    .C(\mem_rdata_latched[29] ),
    .X(_12689_));
 sky130_fd_sc_hd__or3_1 _15364_ (.A(\mem_rdata_latched[26] ),
    .B(\mem_rdata_latched[25] ),
    .C(_12689_),
    .X(_12690_));
 sky130_fd_sc_hd__nor3_2 _15365_ (.A(\mem_rdata_latched[27] ),
    .B(_12688_),
    .C(_12690_),
    .Y(_12691_));
 sky130_vsdinv _15366_ (.A(_12680_),
    .Y(_12692_));
 sky130_fd_sc_hd__o21bai_1 _15367_ (.A1(\mem_rdata_latched[19] ),
    .A2(_12691_),
    .B1_N(_12692_),
    .Y(_12693_));
 sky130_fd_sc_hd__or4_4 _15368_ (.A(\mem_rdata_latched[27] ),
    .B(\mem_rdata_latched[25] ),
    .C(_12689_),
    .D(_12688_),
    .X(_12694_));
 sky130_fd_sc_hd__nand3b_4 _15369_ (.A_N(_12694_),
    .B(\mem_rdata_latched[26] ),
    .C(_12681_),
    .Y(_12695_));
 sky130_fd_sc_hd__o211ai_1 _15370_ (.A1(_00366_),
    .A2(_15210_),
    .B1(_12693_),
    .C1(_12695_),
    .Y(_04066_));
 sky130_vsdinv _15371_ (.A(instr_waitirq),
    .Y(_12696_));
 sky130_fd_sc_hd__nor2_2 _15372_ (.A(decoder_trigger),
    .B(do_waitirq),
    .Y(_12697_));
 sky130_fd_sc_hd__nor2_4 _15373_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .Y(_12698_));
 sky130_fd_sc_hd__and2_1 _15374_ (.A(\cpu_state[1] ),
    .B(decoder_trigger),
    .X(_12699_));
 sky130_vsdinv _15375_ (.A(\irq_pending[31] ),
    .Y(_12700_));
 sky130_vsdinv _15376_ (.A(\irq_mask[29] ),
    .Y(_12701_));
 sky130_fd_sc_hd__nand2_2 _15377_ (.A(_12701_),
    .B(\irq_pending[29] ),
    .Y(_12702_));
 sky130_vsdinv _15378_ (.A(\irq_mask[30] ),
    .Y(_12703_));
 sky130_fd_sc_hd__nand2_2 _15379_ (.A(_12703_),
    .B(\irq_pending[30] ),
    .Y(_12704_));
 sky130_vsdinv _15380_ (.A(\irq_mask[28] ),
    .Y(_12705_));
 sky130_fd_sc_hd__nand2_4 _15381_ (.A(_12705_),
    .B(\irq_pending[28] ),
    .Y(_12706_));
 sky130_fd_sc_hd__o2111ai_4 _15382_ (.A1(\irq_mask[31] ),
    .A2(_12700_),
    .B1(_12702_),
    .C1(_12704_),
    .D1(_12706_),
    .Y(_12707_));
 sky130_vsdinv _15383_ (.A(\irq_pending[14] ),
    .Y(_12708_));
 sky130_vsdinv _15384_ (.A(\irq_mask[12] ),
    .Y(_12709_));
 sky130_fd_sc_hd__nand2_1 _15385_ (.A(_12709_),
    .B(\irq_pending[12] ),
    .Y(_12710_));
 sky130_vsdinv _15386_ (.A(\irq_mask[15] ),
    .Y(_12711_));
 sky130_fd_sc_hd__nand2_4 _15387_ (.A(_12711_),
    .B(\irq_pending[15] ),
    .Y(_12712_));
 sky130_vsdinv _15388_ (.A(\irq_mask[13] ),
    .Y(_12713_));
 sky130_fd_sc_hd__nand2_4 _15389_ (.A(_12713_),
    .B(\irq_pending[13] ),
    .Y(_12714_));
 sky130_fd_sc_hd__o2111ai_4 _15390_ (.A1(\irq_mask[14] ),
    .A2(_12708_),
    .B1(_12710_),
    .C1(_12712_),
    .D1(_12714_),
    .Y(_12715_));
 sky130_fd_sc_hd__nor2_1 _15391_ (.A(_12707_),
    .B(_12715_),
    .Y(_12716_));
 sky130_vsdinv _15392_ (.A(\irq_pending[10] ),
    .Y(_12717_));
 sky130_vsdinv _15393_ (.A(\irq_mask[8] ),
    .Y(_12718_));
 sky130_fd_sc_hd__nand2_1 _15394_ (.A(_12718_),
    .B(\irq_pending[8] ),
    .Y(_12719_));
 sky130_vsdinv _15395_ (.A(\irq_mask[11] ),
    .Y(_12720_));
 sky130_fd_sc_hd__nand2_4 _15396_ (.A(_12720_),
    .B(\irq_pending[11] ),
    .Y(_12721_));
 sky130_vsdinv _15397_ (.A(\irq_mask[9] ),
    .Y(_12722_));
 sky130_fd_sc_hd__nand2_4 _15398_ (.A(_12722_),
    .B(\irq_pending[9] ),
    .Y(_12723_));
 sky130_fd_sc_hd__o2111ai_4 _15399_ (.A1(\irq_mask[10] ),
    .A2(_12717_),
    .B1(_12719_),
    .C1(_12721_),
    .D1(_12723_),
    .Y(_12724_));
 sky130_vsdinv _15400_ (.A(\irq_pending[23] ),
    .Y(_12725_));
 sky130_vsdinv _15401_ (.A(\irq_mask[21] ),
    .Y(_12726_));
 sky130_fd_sc_hd__nand2_2 _15402_ (.A(_12726_),
    .B(\irq_pending[21] ),
    .Y(_12727_));
 sky130_vsdinv _15403_ (.A(\irq_mask[22] ),
    .Y(_12728_));
 sky130_fd_sc_hd__nand2_1 _15404_ (.A(_12728_),
    .B(\irq_pending[22] ),
    .Y(_12729_));
 sky130_vsdinv _15405_ (.A(\irq_mask[20] ),
    .Y(_12730_));
 sky130_fd_sc_hd__nand2_4 _15406_ (.A(_12730_),
    .B(\irq_pending[20] ),
    .Y(_12731_));
 sky130_fd_sc_hd__o2111ai_4 _15407_ (.A1(\irq_mask[23] ),
    .A2(_12725_),
    .B1(_12727_),
    .C1(_12729_),
    .D1(_12731_),
    .Y(_12732_));
 sky130_fd_sc_hd__nor2_1 _15408_ (.A(_12724_),
    .B(_12732_),
    .Y(_12733_));
 sky130_fd_sc_hd__nand2_2 _15409_ (.A(_12716_),
    .B(_12733_),
    .Y(_12734_));
 sky130_vsdinv _15410_ (.A(\irq_pending[6] ),
    .Y(_12735_));
 sky130_vsdinv _15411_ (.A(\irq_mask[4] ),
    .Y(_12736_));
 sky130_fd_sc_hd__nand2_4 _15412_ (.A(_12736_),
    .B(\irq_pending[4] ),
    .Y(_12737_));
 sky130_vsdinv _15413_ (.A(\irq_mask[7] ),
    .Y(_12738_));
 sky130_fd_sc_hd__nand2_4 _15414_ (.A(_12738_),
    .B(\irq_pending[7] ),
    .Y(_12739_));
 sky130_vsdinv _15415_ (.A(\irq_mask[5] ),
    .Y(_12740_));
 sky130_fd_sc_hd__nand2_4 _15416_ (.A(_12740_),
    .B(\irq_pending[5] ),
    .Y(_12741_));
 sky130_fd_sc_hd__o2111ai_4 _15417_ (.A1(\irq_mask[6] ),
    .A2(_12735_),
    .B1(_12737_),
    .C1(_12739_),
    .D1(_12741_),
    .Y(_12742_));
 sky130_vsdinv _15418_ (.A(\irq_pending[27] ),
    .Y(_12743_));
 sky130_vsdinv _15419_ (.A(\irq_mask[25] ),
    .Y(_12744_));
 sky130_fd_sc_hd__nand2_2 _15420_ (.A(_12744_),
    .B(\irq_pending[25] ),
    .Y(_12745_));
 sky130_vsdinv _15421_ (.A(\irq_mask[26] ),
    .Y(_12746_));
 sky130_fd_sc_hd__nand2_4 _15422_ (.A(_12746_),
    .B(\irq_pending[26] ),
    .Y(_12747_));
 sky130_vsdinv _15423_ (.A(\irq_mask[24] ),
    .Y(_12748_));
 sky130_fd_sc_hd__nand2_4 _15424_ (.A(_12748_),
    .B(\irq_pending[24] ),
    .Y(_12749_));
 sky130_fd_sc_hd__o2111ai_4 _15425_ (.A1(\irq_mask[27] ),
    .A2(_12743_),
    .B1(_12745_),
    .C1(_12747_),
    .D1(_12749_),
    .Y(_12750_));
 sky130_fd_sc_hd__nor2_2 _15426_ (.A(_12742_),
    .B(_12750_),
    .Y(_12751_));
 sky130_vsdinv _15427_ (.A(\irq_mask[3] ),
    .Y(_12752_));
 sky130_vsdinv _15428_ (.A(\irq_mask[2] ),
    .Y(_12753_));
 sky130_vsdinv _15429_ (.A(\irq_mask[0] ),
    .Y(_12754_));
 sky130_fd_sc_hd__nand2_2 _15430_ (.A(_12754_),
    .B(\irq_pending[0] ),
    .Y(_12755_));
 sky130_vsdinv _15431_ (.A(\irq_mask[1] ),
    .Y(_12756_));
 sky130_fd_sc_hd__nand2_2 _15432_ (.A(_12756_),
    .B(\irq_pending[1] ),
    .Y(_12757_));
 sky130_fd_sc_hd__nand2_1 _15433_ (.A(_12755_),
    .B(_12757_),
    .Y(_12758_));
 sky130_fd_sc_hd__a221oi_2 _15434_ (.A1(_12752_),
    .A2(\irq_pending[3] ),
    .B1(_12753_),
    .B2(\irq_pending[2] ),
    .C1(_12758_),
    .Y(_12759_));
 sky130_vsdinv _15435_ (.A(\irq_pending[18] ),
    .Y(_12760_));
 sky130_vsdinv _15436_ (.A(\irq_mask[16] ),
    .Y(_12761_));
 sky130_fd_sc_hd__nand2_1 _15437_ (.A(_12761_),
    .B(\irq_pending[16] ),
    .Y(_12762_));
 sky130_vsdinv _15438_ (.A(\irq_mask[19] ),
    .Y(_12763_));
 sky130_fd_sc_hd__nand2_4 _15439_ (.A(_12763_),
    .B(\irq_pending[19] ),
    .Y(_12764_));
 sky130_vsdinv _15440_ (.A(\irq_mask[17] ),
    .Y(_12765_));
 sky130_fd_sc_hd__nand2_2 _15441_ (.A(_12765_),
    .B(\irq_pending[17] ),
    .Y(_12766_));
 sky130_fd_sc_hd__o2111a_1 _15442_ (.A1(\irq_mask[18] ),
    .A2(_12760_),
    .B1(_12762_),
    .C1(_12764_),
    .D1(_12766_),
    .X(_12767_));
 sky130_fd_sc_hd__nand3_4 _15443_ (.A(_12751_),
    .B(_12759_),
    .C(_12767_),
    .Y(_12768_));
 sky130_fd_sc_hd__nor3b_4 _15444_ (.A(irq_active),
    .B(irq_delay),
    .C_N(decoder_trigger),
    .Y(_12769_));
 sky130_vsdinv _15445_ (.A(_12769_),
    .Y(_12770_));
 sky130_fd_sc_hd__o21bai_4 _15446_ (.A1(_12734_),
    .A2(_12768_),
    .B1_N(_12770_),
    .Y(_12771_));
 sky130_fd_sc_hd__o2111ai_4 _15447_ (.A1(_12696_),
    .A2(_12697_),
    .B1(_12698_),
    .C1(_12699_),
    .D1(_12771_),
    .Y(_12772_));
 sky130_vsdinv _15448_ (.A(_12772_),
    .Y(_12773_));
 sky130_fd_sc_hd__o21a_4 _15449_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1(instr_waitirq),
    .X(_00309_));
 sky130_fd_sc_hd__and2_2 _15450_ (.A(_12771_),
    .B(_12698_),
    .X(_12774_));
 sky130_vsdinv _15451_ (.A(_12774_),
    .Y(_00308_));
 sky130_fd_sc_hd__or4b_4 _15452_ (.A(irq_active),
    .B(_00309_),
    .C(_00308_),
    .D_N(_12699_),
    .X(_12775_));
 sky130_fd_sc_hd__o211a_1 _15453_ (.A1(irq_delay),
    .A2(_12773_),
    .B1(_12656_),
    .C1(_12775_),
    .X(_04065_));
 sky130_fd_sc_hd__clkbuf_8 _15454_ (.A(\pcpi_mul.rs1[32] ),
    .X(_12776_));
 sky130_fd_sc_hd__clkbuf_4 _15455_ (.A(_12776_),
    .X(_12777_));
 sky130_fd_sc_hd__buf_6 _15456_ (.A(_12777_),
    .X(_12778_));
 sky130_fd_sc_hd__buf_8 _15457_ (.A(_12778_),
    .X(_12779_));
 sky130_fd_sc_hd__buf_6 _15458_ (.A(_12779_),
    .X(_12780_));
 sky130_fd_sc_hd__buf_4 _15459_ (.A(_12780_),
    .X(_12781_));
 sky130_vsdinv _15460_ (.A(_12781_),
    .Y(_12782_));
 sky130_fd_sc_hd__nor3_4 _15461_ (.A(net293),
    .B(net292),
    .C(net279),
    .Y(_12783_));
 sky130_fd_sc_hd__nand2_1 _15462_ (.A(_12783_),
    .B(net291),
    .Y(_12784_));
 sky130_fd_sc_hd__or3b_2 _15463_ (.A(net296),
    .B(_12784_),
    .C_N(net285),
    .X(_12785_));
 sky130_fd_sc_hd__nor3b_2 _15464_ (.A(net302),
    .B(net299),
    .C_N(net300),
    .Y(_12786_));
 sky130_fd_sc_hd__nand3b_1 _15465_ (.A_N(_12785_),
    .B(net301),
    .C(_12786_),
    .Y(_12787_));
 sky130_fd_sc_hd__nor3_1 _15466_ (.A(net298),
    .B(net297),
    .C(net295),
    .Y(_12788_));
 sky130_fd_sc_hd__and2_2 _15467_ (.A(net101),
    .B(net370),
    .X(_12789_));
 sky130_fd_sc_hd__and3b_2 _15468_ (.A_N(net294),
    .B(_12788_),
    .C(_12789_),
    .X(_12790_));
 sky130_fd_sc_hd__nand3b_4 _15469_ (.A_N(_12787_),
    .B(net274),
    .C(_12790_),
    .Y(_12791_));
 sky130_fd_sc_hd__nor3_4 _15470_ (.A(\pcpi_mul.active[0] ),
    .B(\pcpi_mul.active[1] ),
    .C(_12791_),
    .Y(_12792_));
 sky130_fd_sc_hd__clkbuf_2 _15471_ (.A(_12792_),
    .X(_12793_));
 sky130_fd_sc_hd__clkbuf_4 _15472_ (.A(_12793_),
    .X(_12794_));
 sky130_fd_sc_hd__clkbuf_2 _15473_ (.A(_12792_),
    .X(_12795_));
 sky130_fd_sc_hd__clkbuf_4 _15474_ (.A(_12795_),
    .X(_12796_));
 sky130_fd_sc_hd__clkbuf_4 _15475_ (.A(net330),
    .X(_12797_));
 sky130_fd_sc_hd__nand2_1 _15476_ (.A(_12796_),
    .B(_12797_),
    .Y(_12798_));
 sky130_vsdinv _15477_ (.A(net278),
    .Y(_12799_));
 sky130_fd_sc_hd__nor3_4 _15478_ (.A(_12799_),
    .B(net277),
    .C(_12791_),
    .Y(_12800_));
 sky130_vsdinv _15479_ (.A(net277),
    .Y(_12801_));
 sky130_fd_sc_hd__nor3_4 _15480_ (.A(net278),
    .B(_12801_),
    .C(_12791_),
    .Y(_12802_));
 sky130_fd_sc_hd__nor2_2 _15481_ (.A(_12800_),
    .B(_12802_),
    .Y(_12803_));
 sky130_fd_sc_hd__o22ai_1 _15482_ (.A1(_12782_),
    .A2(_12794_),
    .B1(_12798_),
    .B2(_12803_),
    .Y(_04064_));
 sky130_fd_sc_hd__buf_2 _15483_ (.A(\pcpi_mul.rs2[32] ),
    .X(_12804_));
 sky130_fd_sc_hd__clkbuf_2 _15484_ (.A(_12804_),
    .X(_12805_));
 sky130_vsdinv _15485_ (.A(_12805_),
    .Y(_12806_));
 sky130_fd_sc_hd__buf_1 _15486_ (.A(_12792_),
    .X(_12807_));
 sky130_fd_sc_hd__clkbuf_2 _15487_ (.A(_12807_),
    .X(_03728_));
 sky130_fd_sc_hd__buf_4 _15488_ (.A(net362),
    .X(_12808_));
 sky130_fd_sc_hd__nand3_1 _15489_ (.A(_12802_),
    .B(_12796_),
    .C(_12808_),
    .Y(_12809_));
 sky130_fd_sc_hd__o21ai_1 _15490_ (.A1(_12806_),
    .A2(_03728_),
    .B1(_12809_),
    .Y(_04063_));
 sky130_vsdinv _15491_ (.A(\cpu_state[4] ),
    .Y(_12810_));
 sky130_fd_sc_hd__buf_2 _15492_ (.A(_12810_),
    .X(_12811_));
 sky130_fd_sc_hd__clkbuf_4 _15493_ (.A(_12811_),
    .X(_12812_));
 sky130_fd_sc_hd__buf_2 _15494_ (.A(_12812_),
    .X(_12813_));
 sky130_fd_sc_hd__clkbuf_4 _15495_ (.A(_12643_),
    .X(_12814_));
 sky130_fd_sc_hd__buf_4 _15496_ (.A(_12814_),
    .X(_12815_));
 sky130_fd_sc_hd__and2b_1 _15497_ (.A_N(alu_wait),
    .B(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_12816_));
 sky130_vsdinv _15498_ (.A(_12816_),
    .Y(_12817_));
 sky130_fd_sc_hd__a21oi_1 _15499_ (.A1(_12817_),
    .A2(_00333_),
    .B1(latched_stalu),
    .Y(_12818_));
 sky130_fd_sc_hd__a211oi_1 _15500_ (.A1(_12813_),
    .A2(_00333_),
    .B1(_12815_),
    .C1(_12818_),
    .Y(_04062_));
 sky130_vsdinv _15501_ (.A(\pcpi_mul.active[1] ),
    .Y(_12819_));
 sky130_fd_sc_hd__nor2_4 _15502_ (.A(instr_auipc),
    .B(instr_lui),
    .Y(_12820_));
 sky130_vsdinv _15503_ (.A(instr_jal),
    .Y(_12821_));
 sky130_fd_sc_hd__nand2_2 _15504_ (.A(_12820_),
    .B(_12821_),
    .Y(_00005_));
 sky130_fd_sc_hd__or4_4 _15505_ (.A(instr_lw),
    .B(instr_lh),
    .C(instr_lb),
    .D(instr_jalr),
    .X(_12822_));
 sky130_fd_sc_hd__or4_4 _15506_ (.A(instr_sh),
    .B(instr_sb),
    .C(instr_lhu),
    .D(instr_lbu),
    .X(_12823_));
 sky130_fd_sc_hd__nor3_4 _15507_ (.A(_00005_),
    .B(_12822_),
    .C(_12823_),
    .Y(_12824_));
 sky130_fd_sc_hd__nor2_1 _15508_ (.A(instr_sra),
    .B(instr_srai),
    .Y(_12825_));
 sky130_vsdinv _15509_ (.A(instr_srl),
    .Y(_12826_));
 sky130_vsdinv _15510_ (.A(instr_srli),
    .Y(_12827_));
 sky130_fd_sc_hd__and3_4 _15511_ (.A(_12825_),
    .B(_12826_),
    .C(_12827_),
    .X(_12828_));
 sky130_fd_sc_hd__nand2_8 _15512_ (.A(_12824_),
    .B(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__nor2_8 _15513_ (.A(instr_setq),
    .B(instr_getq),
    .Y(_12830_));
 sky130_vsdinv _15514_ (.A(instr_retirq),
    .Y(_12831_));
 sky130_fd_sc_hd__nand3b_4 _15515_ (.A_N(instr_maskirq),
    .B(_12830_),
    .C(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__or4_4 _15516_ (.A(instr_slt),
    .B(instr_sll),
    .C(instr_sub),
    .D(instr_add),
    .X(_12833_));
 sky130_fd_sc_hd__or4_4 _15517_ (.A(instr_and),
    .B(instr_or),
    .C(instr_xor),
    .D(instr_sltu),
    .X(_12834_));
 sky130_fd_sc_hd__nor3_4 _15518_ (.A(_12832_),
    .B(_12833_),
    .C(_12834_),
    .Y(_12835_));
 sky130_fd_sc_hd__nor3_4 _15519_ (.A(instr_rdinstrh),
    .B(instr_rdinstr),
    .C(instr_rdcycleh),
    .Y(_01714_));
 sky130_fd_sc_hd__nand3b_4 _15520_ (.A_N(instr_rdcycle),
    .B(_12835_),
    .C(net486),
    .Y(_12836_));
 sky130_fd_sc_hd__or4_4 _15521_ (.A(instr_timer),
    .B(instr_waitirq),
    .C(instr_slli),
    .D(instr_sw),
    .X(_12837_));
 sky130_fd_sc_hd__or4_4 _15522_ (.A(instr_slti),
    .B(instr_addi),
    .C(instr_bgeu),
    .D(instr_bltu),
    .X(_12838_));
 sky130_fd_sc_hd__or4_4 _15523_ (.A(instr_andi),
    .B(instr_ori),
    .C(instr_xori),
    .D(instr_sltiu),
    .X(_12839_));
 sky130_fd_sc_hd__or4_4 _15524_ (.A(instr_bge),
    .B(instr_blt),
    .C(instr_bne),
    .D(instr_beq),
    .X(_12840_));
 sky130_fd_sc_hd__or4_4 _15525_ (.A(_12837_),
    .B(_12838_),
    .C(_12839_),
    .D(_12840_),
    .X(_12841_));
 sky130_fd_sc_hd__buf_2 _15526_ (.A(\cpu_state[3] ),
    .X(_12842_));
 sky130_fd_sc_hd__buf_2 _15527_ (.A(_12842_),
    .X(_12843_));
 sky130_fd_sc_hd__o41ai_4 _15528_ (.A1(_12819_),
    .A2(_12829_),
    .A3(_12836_),
    .A4(_12841_),
    .B1(_12843_),
    .Y(_12844_));
 sky130_fd_sc_hd__buf_4 _15529_ (.A(\cpu_state[4] ),
    .X(_12845_));
 sky130_fd_sc_hd__buf_2 _15530_ (.A(alu_wait),
    .X(_12846_));
 sky130_vsdinv _15531_ (.A(\cpu_state[1] ),
    .Y(_12847_));
 sky130_fd_sc_hd__buf_4 _15532_ (.A(_12847_),
    .X(_12848_));
 sky130_fd_sc_hd__clkbuf_4 _15533_ (.A(\cpu_state[2] ),
    .X(_12849_));
 sky130_fd_sc_hd__nor2_2 _15534_ (.A(_12849_),
    .B(\cpu_state[3] ),
    .Y(_12850_));
 sky130_fd_sc_hd__and3_1 _15535_ (.A(_12850_),
    .B(_12810_),
    .C(_12658_),
    .X(_12851_));
 sky130_fd_sc_hd__clkbuf_8 _15536_ (.A(_12851_),
    .X(_01706_));
 sky130_vsdinv _15537_ (.A(_12849_),
    .Y(_12852_));
 sky130_fd_sc_hd__buf_2 _15538_ (.A(_12852_),
    .X(_12853_));
 sky130_fd_sc_hd__or2b_4 _15539_ (.A(instr_rdcycle),
    .B_N(net486),
    .X(_12854_));
 sky130_fd_sc_hd__nor2_8 _15540_ (.A(net494),
    .B(_12832_),
    .Y(_01717_));
 sky130_fd_sc_hd__nor3b_4 _15541_ (.A(_12853_),
    .B(_12854_),
    .C_N(net446),
    .Y(_12855_));
 sky130_fd_sc_hd__a221oi_2 _15542_ (.A1(_12845_),
    .A2(_12846_),
    .B1(_12848_),
    .B2(_01706_),
    .C1(_12855_),
    .Y(_12856_));
 sky130_fd_sc_hd__buf_2 _15543_ (.A(latched_store),
    .X(_12857_));
 sky130_fd_sc_hd__buf_6 _15544_ (.A(_12857_),
    .X(_12858_));
 sky130_fd_sc_hd__a21oi_2 _15545_ (.A1(_12844_),
    .A2(_12856_),
    .B1(_12858_),
    .Y(_12859_));
 sky130_fd_sc_hd__nand3b_1 _15546_ (.A_N(_15244_),
    .B(_12844_),
    .C(_12856_),
    .Y(_12860_));
 sky130_fd_sc_hd__nor3b_4 _15547_ (.A(_12815_),
    .B(_12859_),
    .C_N(_12860_),
    .Y(_04061_));
 sky130_fd_sc_hd__clkbuf_2 _15548_ (.A(\irq_state[1] ),
    .X(_12861_));
 sky130_fd_sc_hd__buf_2 _15549_ (.A(_12861_),
    .X(_12862_));
 sky130_fd_sc_hd__clkbuf_4 _15550_ (.A(\irq_state[0] ),
    .X(_12863_));
 sky130_fd_sc_hd__clkbuf_4 _15551_ (.A(_12863_),
    .X(_12864_));
 sky130_fd_sc_hd__buf_4 _15552_ (.A(\cpu_state[1] ),
    .X(_12865_));
 sky130_fd_sc_hd__buf_4 _15553_ (.A(_12865_),
    .X(_12866_));
 sky130_fd_sc_hd__nand3b_1 _15554_ (.A_N(_12862_),
    .B(_12864_),
    .C(_12866_),
    .Y(_12867_));
 sky130_fd_sc_hd__clkbuf_4 _15555_ (.A(_12848_),
    .X(_12868_));
 sky130_fd_sc_hd__nand2_1 _15556_ (.A(_12868_),
    .B(_12862_),
    .Y(_12869_));
 sky130_fd_sc_hd__clkbuf_4 _15557_ (.A(_12642_),
    .X(_12870_));
 sky130_fd_sc_hd__buf_6 _15558_ (.A(_12870_),
    .X(_12871_));
 sky130_fd_sc_hd__buf_6 _15559_ (.A(_12871_),
    .X(_12872_));
 sky130_fd_sc_hd__a21oi_1 _15560_ (.A1(_12867_),
    .A2(_12869_),
    .B1(_12872_),
    .Y(_04060_));
 sky130_fd_sc_hd__clkbuf_4 _15561_ (.A(_12698_),
    .X(_12873_));
 sky130_fd_sc_hd__o211ai_1 _15562_ (.A1(_12734_),
    .A2(_12768_),
    .B1(_12873_),
    .C1(_12769_),
    .Y(_12874_));
 sky130_fd_sc_hd__buf_4 _15563_ (.A(\cpu_state[1] ),
    .X(_12875_));
 sky130_fd_sc_hd__clkbuf_2 _15564_ (.A(_12875_),
    .X(_12876_));
 sky130_fd_sc_hd__clkbuf_4 _15565_ (.A(_12876_),
    .X(_12877_));
 sky130_fd_sc_hd__buf_2 _15566_ (.A(_12863_),
    .X(_12878_));
 sky130_fd_sc_hd__buf_2 _15567_ (.A(_12865_),
    .X(_12879_));
 sky130_fd_sc_hd__nor2_1 _15568_ (.A(_12878_),
    .B(_12879_),
    .Y(_12880_));
 sky130_fd_sc_hd__a211oi_1 _15569_ (.A1(_12874_),
    .A2(_12877_),
    .B1(_12815_),
    .C1(_12880_),
    .Y(_04059_));
 sky130_fd_sc_hd__o31a_1 _15570_ (.A1(_12829_),
    .A2(_12836_),
    .A3(_12841_),
    .B1(is_lb_lh_lw_lbu_lhu),
    .X(_12881_));
 sky130_fd_sc_hd__nand3_2 _15571_ (.A(_12850_),
    .B(_12810_),
    .C(_12847_),
    .Y(_12882_));
 sky130_fd_sc_hd__o221a_1 _15572_ (.A1(_12811_),
    .A2(_12846_),
    .B1(_12853_),
    .B2(_12881_),
    .C1(_12882_),
    .X(_12883_));
 sky130_vsdinv _15573_ (.A(is_sb_sh_sw),
    .Y(_12884_));
 sky130_fd_sc_hd__nor3_4 _15574_ (.A(_12829_),
    .B(_12836_),
    .C(_12841_),
    .Y(_00310_));
 sky130_fd_sc_hd__clkbuf_4 _15575_ (.A(_12842_),
    .X(_12885_));
 sky130_fd_sc_hd__nor2_4 _15576_ (.A(_12829_),
    .B(_12841_),
    .Y(_12886_));
 sky130_fd_sc_hd__and2b_1 _15577_ (.A_N(_12854_),
    .B(_12835_),
    .X(_12887_));
 sky130_fd_sc_hd__nand3_1 _15578_ (.A(_12886_),
    .B(\pcpi_mul.active[1] ),
    .C(_12887_),
    .Y(_12888_));
 sky130_fd_sc_hd__o211ai_2 _15579_ (.A1(_12884_),
    .A2(_00310_),
    .B1(_12885_),
    .C1(_12888_),
    .Y(_12889_));
 sky130_fd_sc_hd__a21oi_4 _15580_ (.A1(_12632_),
    .A2(net456),
    .B1(_12641_),
    .Y(_12890_));
 sky130_vsdinv _15581_ (.A(_12890_),
    .Y(_12891_));
 sky130_fd_sc_hd__a21oi_2 _15582_ (.A1(_12883_),
    .A2(_12889_),
    .B1(_12891_),
    .Y(_12892_));
 sky130_vsdinv _15583_ (.A(\cpu_state[0] ),
    .Y(_12893_));
 sky130_fd_sc_hd__and3_1 _15584_ (.A(_12850_),
    .B(_12847_),
    .C(_12893_),
    .X(_12894_));
 sky130_fd_sc_hd__buf_2 _15585_ (.A(_12648_),
    .X(_12895_));
 sky130_vsdinv _15586_ (.A(_00343_),
    .Y(_12896_));
 sky130_fd_sc_hd__nor2_8 _15587_ (.A(\cpu_state[6] ),
    .B(\cpu_state[5] ),
    .Y(_00297_));
 sky130_fd_sc_hd__and4_1 _15588_ (.A(_12816_),
    .B(_12895_),
    .C(_12896_),
    .D(_00297_),
    .X(_12897_));
 sky130_fd_sc_hd__nor3_2 _15589_ (.A(_00356_),
    .B(_12891_),
    .C(_12892_),
    .Y(_12898_));
 sky130_fd_sc_hd__a221o_1 _15590_ (.A1(_12666_),
    .A2(_12892_),
    .B1(_12894_),
    .B2(_12897_),
    .C1(_12898_),
    .X(_04058_));
 sky130_fd_sc_hd__buf_2 _15591_ (.A(instr_jal),
    .X(_12899_));
 sky130_fd_sc_hd__clkbuf_4 _15592_ (.A(_12899_),
    .X(_12900_));
 sky130_fd_sc_hd__clkbuf_4 _15593_ (.A(_12772_),
    .X(_12901_));
 sky130_fd_sc_hd__nor2_1 _15594_ (.A(_12900_),
    .B(_12901_),
    .Y(_12902_));
 sky130_fd_sc_hd__buf_4 _15595_ (.A(_12821_),
    .X(_00323_));
 sky130_fd_sc_hd__o211ai_2 _15596_ (.A1(instr_retirq),
    .A2(instr_jalr),
    .B1(_00323_),
    .C1(_12773_),
    .Y(_12903_));
 sky130_fd_sc_hd__o211a_1 _15597_ (.A1(_12640_),
    .A2(_12902_),
    .B1(_12890_),
    .C1(_12903_),
    .X(_04057_));
 sky130_fd_sc_hd__nor3b_2 _15598_ (.A(net480),
    .B(net478),
    .C_N(net449),
    .Y(_12904_));
 sky130_fd_sc_hd__nor3b_4 _15599_ (.A(_00358_),
    .B(_00357_),
    .C_N(_12904_),
    .Y(_12905_));
 sky130_fd_sc_hd__buf_2 _15600_ (.A(_12905_),
    .X(_12906_));
 sky130_fd_sc_hd__clkbuf_4 _15601_ (.A(_12906_),
    .X(_12907_));
 sky130_fd_sc_hd__nor2_8 _15602_ (.A(_01207_),
    .B(net425),
    .Y(\cpuregs_rs1[31] ));
 sky130_fd_sc_hd__clkbuf_2 _15603_ (.A(instr_maskirq),
    .X(_12908_));
 sky130_fd_sc_hd__and2_1 _15604_ (.A(_12908_),
    .B(_12849_),
    .X(_12909_));
 sky130_fd_sc_hd__buf_2 _15605_ (.A(_12909_),
    .X(_12910_));
 sky130_fd_sc_hd__clkbuf_2 _15606_ (.A(_12910_),
    .X(_12911_));
 sky130_fd_sc_hd__buf_4 _15607_ (.A(_12642_),
    .X(_12912_));
 sky130_fd_sc_hd__clkbuf_2 _15608_ (.A(_12912_),
    .X(_12913_));
 sky130_fd_sc_hd__buf_2 _15609_ (.A(_12908_),
    .X(_12914_));
 sky130_fd_sc_hd__clkbuf_4 _15610_ (.A(_12849_),
    .X(_12915_));
 sky130_fd_sc_hd__buf_4 _15611_ (.A(_12915_),
    .X(_12916_));
 sky130_fd_sc_hd__clkbuf_4 _15612_ (.A(_12916_),
    .X(_12917_));
 sky130_fd_sc_hd__a21boi_1 _15613_ (.A1(_12914_),
    .A2(_12917_),
    .B1_N(\irq_mask[31] ),
    .Y(_12918_));
 sky130_fd_sc_hd__a211o_1 _15614_ (.A1(\cpuregs_rs1[31] ),
    .A2(_12911_),
    .B1(_12913_),
    .C1(_12918_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_2 _15615_ (.A(_12910_),
    .X(_12919_));
 sky130_fd_sc_hd__buf_4 _15616_ (.A(_12895_),
    .X(_12920_));
 sky130_fd_sc_hd__clkbuf_2 _15617_ (.A(_12920_),
    .X(_12921_));
 sky130_fd_sc_hd__clkbuf_8 _15618_ (.A(_12906_),
    .X(_12922_));
 sky130_fd_sc_hd__nor2_8 _15619_ (.A(_01180_),
    .B(_12922_),
    .Y(\cpuregs_rs1[30] ));
 sky130_fd_sc_hd__clkbuf_2 _15620_ (.A(_12909_),
    .X(_12923_));
 sky130_fd_sc_hd__buf_2 _15621_ (.A(_12923_),
    .X(_12924_));
 sky130_fd_sc_hd__nand2_1 _15622_ (.A(\cpuregs_rs1[30] ),
    .B(_12924_),
    .Y(_12925_));
 sky130_fd_sc_hd__o211ai_1 _15623_ (.A1(_12703_),
    .A2(_12919_),
    .B1(_12921_),
    .C1(_12925_),
    .Y(_04055_));
 sky130_fd_sc_hd__nor2_8 _15624_ (.A(_01153_),
    .B(_12922_),
    .Y(\cpuregs_rs1[29] ));
 sky130_fd_sc_hd__nand2_1 _15625_ (.A(\cpuregs_rs1[29] ),
    .B(_12924_),
    .Y(_12926_));
 sky130_fd_sc_hd__o211ai_1 _15626_ (.A1(_12701_),
    .A2(_12919_),
    .B1(_12921_),
    .C1(_12926_),
    .Y(_04054_));
 sky130_fd_sc_hd__buf_4 _15627_ (.A(_12905_),
    .X(_12927_));
 sky130_fd_sc_hd__nor2_8 _15628_ (.A(_01126_),
    .B(net434),
    .Y(\cpuregs_rs1[28] ));
 sky130_fd_sc_hd__nand2_1 _15629_ (.A(\cpuregs_rs1[28] ),
    .B(_12924_),
    .Y(_12928_));
 sky130_fd_sc_hd__o211ai_1 _15630_ (.A1(_12705_),
    .A2(_12919_),
    .B1(_12921_),
    .C1(_12928_),
    .Y(_04053_));
 sky130_fd_sc_hd__nor2_8 _15631_ (.A(_01099_),
    .B(net425),
    .Y(\cpuregs_rs1[27] ));
 sky130_fd_sc_hd__clkbuf_2 _15632_ (.A(_12916_),
    .X(_12929_));
 sky130_fd_sc_hd__a21boi_1 _15633_ (.A1(_12914_),
    .A2(_12929_),
    .B1_N(\irq_mask[27] ),
    .Y(_12930_));
 sky130_fd_sc_hd__a211o_1 _15634_ (.A1(\cpuregs_rs1[27] ),
    .A2(_12911_),
    .B1(_12913_),
    .C1(_12930_),
    .X(_04052_));
 sky130_fd_sc_hd__nor2_8 _15635_ (.A(_01072_),
    .B(net434),
    .Y(\cpuregs_rs1[26] ));
 sky130_fd_sc_hd__nand2_1 _15636_ (.A(\cpuregs_rs1[26] ),
    .B(_12924_),
    .Y(_12931_));
 sky130_fd_sc_hd__o211ai_1 _15637_ (.A1(_12746_),
    .A2(_12919_),
    .B1(_12921_),
    .C1(_12931_),
    .Y(_04051_));
 sky130_fd_sc_hd__nor2_8 _15638_ (.A(_01045_),
    .B(_12927_),
    .Y(\cpuregs_rs1[25] ));
 sky130_fd_sc_hd__clkbuf_2 _15639_ (.A(_12923_),
    .X(_12932_));
 sky130_fd_sc_hd__nand2_1 _15640_ (.A(\cpuregs_rs1[25] ),
    .B(_12932_),
    .Y(_12933_));
 sky130_fd_sc_hd__o211ai_1 _15641_ (.A1(_12744_),
    .A2(_12919_),
    .B1(_12921_),
    .C1(_12933_),
    .Y(_04050_));
 sky130_fd_sc_hd__nor2_8 _15642_ (.A(_01018_),
    .B(net434),
    .Y(\cpuregs_rs1[24] ));
 sky130_fd_sc_hd__nand2_1 _15643_ (.A(\cpuregs_rs1[24] ),
    .B(_12932_),
    .Y(_12934_));
 sky130_fd_sc_hd__o211ai_1 _15644_ (.A1(_12748_),
    .A2(_12919_),
    .B1(_12921_),
    .C1(_12934_),
    .Y(_04049_));
 sky130_fd_sc_hd__nor2_8 _15645_ (.A(_00991_),
    .B(net425),
    .Y(\cpuregs_rs1[23] ));
 sky130_fd_sc_hd__a21boi_1 _15646_ (.A1(_12914_),
    .A2(_12929_),
    .B1_N(\irq_mask[23] ),
    .Y(_12935_));
 sky130_fd_sc_hd__a211o_1 _15647_ (.A1(\cpuregs_rs1[23] ),
    .A2(_12911_),
    .B1(_12913_),
    .C1(_12935_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_2 _15648_ (.A(_12910_),
    .X(_12936_));
 sky130_fd_sc_hd__clkbuf_2 _15649_ (.A(_12920_),
    .X(_12937_));
 sky130_fd_sc_hd__nor2_8 _15650_ (.A(_00964_),
    .B(_12927_),
    .Y(\cpuregs_rs1[22] ));
 sky130_fd_sc_hd__nand2_1 _15651_ (.A(\cpuregs_rs1[22] ),
    .B(_12932_),
    .Y(_12938_));
 sky130_fd_sc_hd__o211ai_1 _15652_ (.A1(_12728_),
    .A2(_12936_),
    .B1(_12937_),
    .C1(_12938_),
    .Y(_04047_));
 sky130_fd_sc_hd__nor2_8 _15653_ (.A(_00937_),
    .B(net434),
    .Y(\cpuregs_rs1[21] ));
 sky130_fd_sc_hd__nand2_1 _15654_ (.A(\cpuregs_rs1[21] ),
    .B(_12932_),
    .Y(_12939_));
 sky130_fd_sc_hd__o211ai_1 _15655_ (.A1(_12726_),
    .A2(_12936_),
    .B1(_12937_),
    .C1(_12939_),
    .Y(_04046_));
 sky130_fd_sc_hd__buf_6 _15656_ (.A(_12905_),
    .X(_12940_));
 sky130_fd_sc_hd__nor2_8 _15657_ (.A(_00910_),
    .B(_12940_),
    .Y(\cpuregs_rs1[20] ));
 sky130_fd_sc_hd__nand2_1 _15658_ (.A(\cpuregs_rs1[20] ),
    .B(_12932_),
    .Y(_12941_));
 sky130_fd_sc_hd__o211ai_1 _15659_ (.A1(_12730_),
    .A2(_12936_),
    .B1(_12937_),
    .C1(_12941_),
    .Y(_04045_));
 sky130_fd_sc_hd__nor2_8 _15660_ (.A(_00883_),
    .B(net433),
    .Y(\cpuregs_rs1[19] ));
 sky130_fd_sc_hd__nand2_1 _15661_ (.A(\cpuregs_rs1[19] ),
    .B(_12932_),
    .Y(_12942_));
 sky130_fd_sc_hd__o211ai_1 _15662_ (.A1(_12763_),
    .A2(_12936_),
    .B1(_12937_),
    .C1(_12942_),
    .Y(_04044_));
 sky130_fd_sc_hd__nor2_8 _15663_ (.A(_00856_),
    .B(net424),
    .Y(\cpuregs_rs1[18] ));
 sky130_fd_sc_hd__a21boi_1 _15664_ (.A1(_12914_),
    .A2(_12929_),
    .B1_N(\irq_mask[18] ),
    .Y(_12943_));
 sky130_fd_sc_hd__a211o_1 _15665_ (.A1(\cpuregs_rs1[18] ),
    .A2(_12911_),
    .B1(_12913_),
    .C1(_12943_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_8 _15666_ (.A(_00829_),
    .B(_12940_),
    .Y(\cpuregs_rs1[17] ));
 sky130_fd_sc_hd__clkbuf_2 _15667_ (.A(_12923_),
    .X(_12944_));
 sky130_fd_sc_hd__nand2_1 _15668_ (.A(\cpuregs_rs1[17] ),
    .B(_12944_),
    .Y(_12945_));
 sky130_fd_sc_hd__o211ai_1 _15669_ (.A1(_12765_),
    .A2(_12936_),
    .B1(_12937_),
    .C1(_12945_),
    .Y(_04042_));
 sky130_fd_sc_hd__nor2_8 _15670_ (.A(_00802_),
    .B(net433),
    .Y(\cpuregs_rs1[16] ));
 sky130_fd_sc_hd__nand2_1 _15671_ (.A(\cpuregs_rs1[16] ),
    .B(_12944_),
    .Y(_12946_));
 sky130_fd_sc_hd__o211ai_1 _15672_ (.A1(_12761_),
    .A2(_12936_),
    .B1(_12937_),
    .C1(_12946_),
    .Y(_04041_));
 sky130_fd_sc_hd__clkbuf_2 _15673_ (.A(_12923_),
    .X(_12947_));
 sky130_fd_sc_hd__clkbuf_2 _15674_ (.A(_12920_),
    .X(_12948_));
 sky130_fd_sc_hd__nor2_8 _15675_ (.A(_00775_),
    .B(net433),
    .Y(\cpuregs_rs1[15] ));
 sky130_fd_sc_hd__nand2_1 _15676_ (.A(\cpuregs_rs1[15] ),
    .B(_12944_),
    .Y(_12949_));
 sky130_fd_sc_hd__o211ai_1 _15677_ (.A1(_12711_),
    .A2(_12947_),
    .B1(_12948_),
    .C1(_12949_),
    .Y(_04040_));
 sky130_fd_sc_hd__nor2_8 _15678_ (.A(_00748_),
    .B(net424),
    .Y(\cpuregs_rs1[14] ));
 sky130_fd_sc_hd__a21boi_1 _15679_ (.A1(_12914_),
    .A2(_12929_),
    .B1_N(\irq_mask[14] ),
    .Y(_12950_));
 sky130_fd_sc_hd__a211o_1 _15680_ (.A1(\cpuregs_rs1[14] ),
    .A2(_12911_),
    .B1(_12913_),
    .C1(_12950_),
    .X(_04039_));
 sky130_fd_sc_hd__nor2_8 _15681_ (.A(_00721_),
    .B(net433),
    .Y(\cpuregs_rs1[13] ));
 sky130_fd_sc_hd__nand2_1 _15682_ (.A(\cpuregs_rs1[13] ),
    .B(_12944_),
    .Y(_12951_));
 sky130_fd_sc_hd__o211ai_1 _15683_ (.A1(_12713_),
    .A2(_12947_),
    .B1(_12948_),
    .C1(_12951_),
    .Y(_04038_));
 sky130_fd_sc_hd__buf_4 _15684_ (.A(_12905_),
    .X(_12952_));
 sky130_fd_sc_hd__nor2_8 _15685_ (.A(_00694_),
    .B(net432),
    .Y(\cpuregs_rs1[12] ));
 sky130_fd_sc_hd__nand2_1 _15686_ (.A(\cpuregs_rs1[12] ),
    .B(_12944_),
    .Y(_12953_));
 sky130_fd_sc_hd__o211ai_1 _15687_ (.A1(_12709_),
    .A2(_12947_),
    .B1(_12948_),
    .C1(_12953_),
    .Y(_04037_));
 sky130_fd_sc_hd__nor2_8 _15688_ (.A(_00667_),
    .B(net432),
    .Y(\cpuregs_rs1[11] ));
 sky130_fd_sc_hd__nand2_1 _15689_ (.A(\cpuregs_rs1[11] ),
    .B(_12944_),
    .Y(_12954_));
 sky130_fd_sc_hd__o211ai_1 _15690_ (.A1(_12720_),
    .A2(_12947_),
    .B1(_12948_),
    .C1(_12954_),
    .Y(_04036_));
 sky130_fd_sc_hd__nor2_8 _15691_ (.A(_00640_),
    .B(net424),
    .Y(\cpuregs_rs1[10] ));
 sky130_fd_sc_hd__clkbuf_2 _15692_ (.A(_12908_),
    .X(_12955_));
 sky130_fd_sc_hd__a21boi_1 _15693_ (.A1(_12955_),
    .A2(_12929_),
    .B1_N(\irq_mask[10] ),
    .Y(_12956_));
 sky130_fd_sc_hd__a211o_1 _15694_ (.A1(\cpuregs_rs1[10] ),
    .A2(_12924_),
    .B1(_12913_),
    .C1(_12956_),
    .X(_04035_));
 sky130_fd_sc_hd__nor2_8 _15695_ (.A(_00613_),
    .B(_12952_),
    .Y(\cpuregs_rs1[9] ));
 sky130_fd_sc_hd__clkbuf_2 _15696_ (.A(_12923_),
    .X(_12957_));
 sky130_fd_sc_hd__nand2_1 _15697_ (.A(\cpuregs_rs1[9] ),
    .B(_12957_),
    .Y(_12958_));
 sky130_fd_sc_hd__o211ai_1 _15698_ (.A1(_12722_),
    .A2(_12947_),
    .B1(_12948_),
    .C1(_12958_),
    .Y(_04034_));
 sky130_fd_sc_hd__nor2_8 _15699_ (.A(_00586_),
    .B(net432),
    .Y(\cpuregs_rs1[8] ));
 sky130_fd_sc_hd__nand2_1 _15700_ (.A(\cpuregs_rs1[8] ),
    .B(_12957_),
    .Y(_12959_));
 sky130_fd_sc_hd__o211ai_1 _15701_ (.A1(_12718_),
    .A2(_12947_),
    .B1(_12948_),
    .C1(_12959_),
    .Y(_04033_));
 sky130_fd_sc_hd__clkbuf_2 _15702_ (.A(_12923_),
    .X(_12960_));
 sky130_fd_sc_hd__clkbuf_4 _15703_ (.A(_12654_),
    .X(_12961_));
 sky130_fd_sc_hd__clkbuf_2 _15704_ (.A(_12961_),
    .X(_12962_));
 sky130_fd_sc_hd__nor2_8 _15705_ (.A(_00559_),
    .B(_12952_),
    .Y(\cpuregs_rs1[7] ));
 sky130_fd_sc_hd__nand2_1 _15706_ (.A(\cpuregs_rs1[7] ),
    .B(_12957_),
    .Y(_12963_));
 sky130_fd_sc_hd__o211ai_1 _15707_ (.A1(_12738_),
    .A2(_12960_),
    .B1(_12962_),
    .C1(_12963_),
    .Y(_04032_));
 sky130_fd_sc_hd__nor2_8 _15708_ (.A(_00532_),
    .B(net424),
    .Y(\cpuregs_rs1[6] ));
 sky130_fd_sc_hd__buf_6 _15709_ (.A(_12912_),
    .X(_12964_));
 sky130_fd_sc_hd__a21boi_1 _15710_ (.A1(_12955_),
    .A2(_12929_),
    .B1_N(\irq_mask[6] ),
    .Y(_12965_));
 sky130_fd_sc_hd__a211o_1 _15711_ (.A1(\cpuregs_rs1[6] ),
    .A2(_12924_),
    .B1(_12964_),
    .C1(_12965_),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_8 _15712_ (.A(_00505_),
    .B(net432),
    .Y(\cpuregs_rs1[5] ));
 sky130_fd_sc_hd__nand2_1 _15713_ (.A(\cpuregs_rs1[5] ),
    .B(_12957_),
    .Y(_12966_));
 sky130_fd_sc_hd__o211ai_1 _15714_ (.A1(_12740_),
    .A2(_12960_),
    .B1(_12962_),
    .C1(_12966_),
    .Y(_04030_));
 sky130_fd_sc_hd__nor2_8 _15715_ (.A(_00478_),
    .B(net435),
    .Y(\cpuregs_rs1[4] ));
 sky130_fd_sc_hd__nand2_1 _15716_ (.A(\cpuregs_rs1[4] ),
    .B(_12957_),
    .Y(_12967_));
 sky130_fd_sc_hd__o211ai_1 _15717_ (.A1(_12736_),
    .A2(_12960_),
    .B1(_12962_),
    .C1(_12967_),
    .Y(_04029_));
 sky130_fd_sc_hd__nor2_8 _15718_ (.A(_00451_),
    .B(net435),
    .Y(\cpuregs_rs1[3] ));
 sky130_fd_sc_hd__nand2_1 _15719_ (.A(\cpuregs_rs1[3] ),
    .B(_12957_),
    .Y(_12968_));
 sky130_fd_sc_hd__o211ai_1 _15720_ (.A1(_12752_),
    .A2(_12960_),
    .B1(_12962_),
    .C1(_12968_),
    .Y(_04028_));
 sky130_fd_sc_hd__nor2_8 _15721_ (.A(_00424_),
    .B(net435),
    .Y(\cpuregs_rs1[2] ));
 sky130_fd_sc_hd__nand2_1 _15722_ (.A(\cpuregs_rs1[2] ),
    .B(_12910_),
    .Y(_12969_));
 sky130_fd_sc_hd__o211ai_1 _15723_ (.A1(_12753_),
    .A2(_12960_),
    .B1(_12962_),
    .C1(_12969_),
    .Y(_04027_));
 sky130_fd_sc_hd__nor2_8 _15724_ (.A(_00397_),
    .B(net435),
    .Y(\cpuregs_rs1[1] ));
 sky130_fd_sc_hd__nand2_1 _15725_ (.A(\cpuregs_rs1[1] ),
    .B(_12910_),
    .Y(_12970_));
 sky130_fd_sc_hd__o211ai_1 _15726_ (.A1(_12756_),
    .A2(_12960_),
    .B1(_12962_),
    .C1(_12970_),
    .Y(_04026_));
 sky130_fd_sc_hd__buf_2 _15727_ (.A(_12920_),
    .X(_12971_));
 sky130_fd_sc_hd__nand3b_1 _15728_ (.A_N(_12907_),
    .B(_00370_),
    .C(_12910_),
    .Y(_12972_));
 sky130_fd_sc_hd__o211ai_1 _15729_ (.A1(_12754_),
    .A2(_12911_),
    .B1(_12971_),
    .C1(_12972_),
    .Y(_04025_));
 sky130_fd_sc_hd__nor2b_4 _15730_ (.A(_12907_),
    .B_N(_00370_),
    .Y(\cpuregs_rs1[0] ));
 sky130_fd_sc_hd__a21boi_4 _15731_ (.A1(_12635_),
    .A2(_12670_),
    .B1_N(_00290_),
    .Y(_12973_));
 sky130_fd_sc_hd__nand2_8 _15732_ (.A(_12973_),
    .B(_12675_),
    .Y(_12974_));
 sky130_fd_sc_hd__buf_4 _15733_ (.A(_12974_),
    .X(_12975_));
 sky130_fd_sc_hd__clkbuf_4 _15734_ (.A(mem_do_wdata),
    .X(_12976_));
 sky130_fd_sc_hd__clkinv_4 _15735_ (.A(_12976_),
    .Y(_00291_));
 sky130_fd_sc_hd__o2111a_2 _15736_ (.A1(_12666_),
    .A2(_12640_),
    .B1(_00291_),
    .C1(_12675_),
    .D1(_12973_),
    .X(_12977_));
 sky130_fd_sc_hd__a21o_1 _15737_ (.A1(net166),
    .A2(_12975_),
    .B1(_12977_),
    .X(_04024_));
 sky130_fd_sc_hd__buf_2 _15738_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_12978_));
 sky130_fd_sc_hd__buf_2 _15739_ (.A(_12978_),
    .X(_12979_));
 sky130_fd_sc_hd__buf_2 _15740_ (.A(_12979_),
    .X(_12980_));
 sky130_fd_sc_hd__buf_2 _15741_ (.A(_12681_),
    .X(_12981_));
 sky130_fd_sc_hd__nand3b_4 _15742_ (.A_N(_00328_),
    .B(_00329_),
    .C(_00330_),
    .Y(_12982_));
 sky130_fd_sc_hd__o31ai_1 _15743_ (.A1(_00327_),
    .A2(_12683_),
    .A3(_12982_),
    .B1(_12681_),
    .Y(_12983_));
 sky130_fd_sc_hd__o211a_1 _15744_ (.A1(_12980_),
    .A2(_12981_),
    .B1(_12656_),
    .C1(_12983_),
    .X(_04023_));
 sky130_fd_sc_hd__clkbuf_2 _15745_ (.A(_12692_),
    .X(_12984_));
 sky130_fd_sc_hd__buf_4 _15746_ (.A(_12984_),
    .X(_00337_));
 sky130_fd_sc_hd__nand2b_2 _15747_ (.A_N(_12694_),
    .B(\mem_rdata_latched[26] ),
    .Y(_12985_));
 sky130_fd_sc_hd__nand3_1 _15748_ (.A(_12985_),
    .B(\mem_rdata_latched[18] ),
    .C(_12981_),
    .Y(_12986_));
 sky130_fd_sc_hd__a21bo_1 _15749_ (.A1(\decoded_rs1[3] ),
    .A2(_00337_),
    .B1_N(_12986_),
    .X(_04022_));
 sky130_fd_sc_hd__nand3_1 _15750_ (.A(_12985_),
    .B(\mem_rdata_latched[17] ),
    .C(_12981_),
    .Y(_12987_));
 sky130_fd_sc_hd__a21bo_1 _15751_ (.A1(\decoded_rs1[2] ),
    .A2(_00337_),
    .B1_N(_12987_),
    .X(_04021_));
 sky130_fd_sc_hd__nand3_1 _15752_ (.A(_12985_),
    .B(\mem_rdata_latched[16] ),
    .C(_12981_),
    .Y(_12988_));
 sky130_fd_sc_hd__a21bo_1 _15753_ (.A1(\decoded_rs1[1] ),
    .A2(_00337_),
    .B1_N(_12988_),
    .X(_04020_));
 sky130_fd_sc_hd__nand3_1 _15754_ (.A(_12985_),
    .B(\mem_rdata_latched[15] ),
    .C(_12981_),
    .Y(_12989_));
 sky130_fd_sc_hd__a21bo_1 _15755_ (.A1(\decoded_rs1[0] ),
    .A2(_00337_),
    .B1_N(_12989_),
    .X(_04019_));
 sky130_fd_sc_hd__clkbuf_4 _15756_ (.A(\mem_rdata_q[14] ),
    .X(_12990_));
 sky130_fd_sc_hd__clkbuf_4 _15757_ (.A(\mem_rdata_q[13] ),
    .X(_12991_));
 sky130_fd_sc_hd__clkbuf_4 _15758_ (.A(_12991_),
    .X(_12992_));
 sky130_fd_sc_hd__buf_2 _15759_ (.A(\mem_rdata_q[12] ),
    .X(_12993_));
 sky130_fd_sc_hd__clkbuf_4 _15760_ (.A(_12993_),
    .X(_12994_));
 sky130_fd_sc_hd__nand3_2 _15761_ (.A(_12990_),
    .B(_12992_),
    .C(_12994_),
    .Y(_12995_));
 sky130_fd_sc_hd__nor3_4 _15762_ (.A(\mem_rdata_q[31] ),
    .B(\mem_rdata_q[30] ),
    .C(\mem_rdata_q[29] ),
    .Y(_12996_));
 sky130_fd_sc_hd__clkbuf_4 _15763_ (.A(decoder_trigger),
    .X(_12997_));
 sky130_fd_sc_hd__and2b_1 _15764_ (.A_N(decoder_pseudo_trigger),
    .B(_12997_),
    .X(_12998_));
 sky130_fd_sc_hd__nor2_2 _15765_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[26] ),
    .Y(_12999_));
 sky130_fd_sc_hd__nor2_2 _15766_ (.A(\mem_rdata_q[27] ),
    .B(\mem_rdata_q[25] ),
    .Y(_13000_));
 sky130_fd_sc_hd__and4_1 _15767_ (.A(_12996_),
    .B(_12998_),
    .C(_12999_),
    .D(_13000_),
    .X(_13001_));
 sky130_fd_sc_hd__clkbuf_2 _15768_ (.A(_13001_),
    .X(_13002_));
 sky130_fd_sc_hd__nand3b_1 _15769_ (.A_N(_12995_),
    .B(_13002_),
    .C(is_alu_reg_reg),
    .Y(_13003_));
 sky130_vsdinv _15770_ (.A(_12998_),
    .Y(_13004_));
 sky130_fd_sc_hd__clkbuf_4 _15771_ (.A(_13004_),
    .X(_13005_));
 sky130_fd_sc_hd__clkbuf_2 _15772_ (.A(_13005_),
    .X(_13006_));
 sky130_fd_sc_hd__clkbuf_4 _15773_ (.A(instr_and),
    .X(_13007_));
 sky130_fd_sc_hd__nand2_1 _15774_ (.A(_13006_),
    .B(_13007_),
    .Y(_13008_));
 sky130_fd_sc_hd__clkbuf_2 _15775_ (.A(_12871_),
    .X(_13009_));
 sky130_fd_sc_hd__a21oi_1 _15776_ (.A1(_13003_),
    .A2(_13008_),
    .B1(_13009_),
    .Y(_04018_));
 sky130_fd_sc_hd__nand3b_4 _15777_ (.A_N(_12993_),
    .B(_12990_),
    .C(_12991_),
    .Y(_13010_));
 sky130_fd_sc_hd__nand3b_1 _15778_ (.A_N(_13010_),
    .B(_13002_),
    .C(is_alu_reg_reg),
    .Y(_13011_));
 sky130_fd_sc_hd__buf_4 _15779_ (.A(instr_or),
    .X(_13012_));
 sky130_fd_sc_hd__nand2_1 _15780_ (.A(_13006_),
    .B(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__a21oi_1 _15781_ (.A1(_13011_),
    .A2(_13013_),
    .B1(_13009_),
    .Y(_04017_));
 sky130_fd_sc_hd__clkbuf_4 _15782_ (.A(\mem_rdata_q[29] ),
    .X(_13014_));
 sky130_vsdinv _15783_ (.A(\mem_rdata_q[30] ),
    .Y(_13015_));
 sky130_vsdinv _15784_ (.A(_12999_),
    .Y(_13016_));
 sky130_fd_sc_hd__or4b_4 _15785_ (.A(\mem_rdata_q[31] ),
    .B(_13015_),
    .C(_13016_),
    .D_N(_13000_),
    .X(_13017_));
 sky130_fd_sc_hd__nor3_4 _15786_ (.A(_13014_),
    .B(_13005_),
    .C(_13017_),
    .Y(_13018_));
 sky130_fd_sc_hd__buf_2 _15787_ (.A(is_alu_reg_reg),
    .X(_13019_));
 sky130_fd_sc_hd__nand3b_4 _15788_ (.A_N(_12991_),
    .B(\mem_rdata_q[14] ),
    .C(_12993_),
    .Y(_13020_));
 sky130_vsdinv _15789_ (.A(_13020_),
    .Y(_13021_));
 sky130_fd_sc_hd__nand3_2 _15790_ (.A(_13018_),
    .B(_13019_),
    .C(_13021_),
    .Y(_13022_));
 sky130_fd_sc_hd__nand2_1 _15791_ (.A(_13006_),
    .B(instr_sra),
    .Y(_13023_));
 sky130_fd_sc_hd__a21oi_1 _15792_ (.A1(_13022_),
    .A2(_13023_),
    .B1(_13009_),
    .Y(_04016_));
 sky130_fd_sc_hd__buf_2 _15793_ (.A(_13001_),
    .X(_13024_));
 sky130_fd_sc_hd__nand3_1 _15794_ (.A(_13024_),
    .B(_13019_),
    .C(_13021_),
    .Y(_13025_));
 sky130_fd_sc_hd__nand2_1 _15795_ (.A(_13006_),
    .B(instr_srl),
    .Y(_13026_));
 sky130_fd_sc_hd__a21oi_1 _15796_ (.A1(_13025_),
    .A2(_13026_),
    .B1(_13009_),
    .Y(_04015_));
 sky130_fd_sc_hd__nor3b_4 _15797_ (.A(_12992_),
    .B(_12994_),
    .C_N(_12990_),
    .Y(_13027_));
 sky130_fd_sc_hd__nand3_2 _15798_ (.A(_13024_),
    .B(_13019_),
    .C(_13027_),
    .Y(_13028_));
 sky130_fd_sc_hd__nand2_1 _15799_ (.A(_13006_),
    .B(instr_xor),
    .Y(_13029_));
 sky130_fd_sc_hd__a21oi_1 _15800_ (.A1(_13028_),
    .A2(_13029_),
    .B1(_13009_),
    .Y(_04014_));
 sky130_fd_sc_hd__and3b_1 _15801_ (.A_N(\mem_rdata_q[14] ),
    .B(_12991_),
    .C(_12993_),
    .X(_13030_));
 sky130_fd_sc_hd__nand3_1 _15802_ (.A(_13002_),
    .B(_13019_),
    .C(_13030_),
    .Y(_13031_));
 sky130_fd_sc_hd__nand2_1 _15803_ (.A(_13006_),
    .B(instr_sltu),
    .Y(_13032_));
 sky130_fd_sc_hd__a21oi_1 _15804_ (.A1(_13031_),
    .A2(_13032_),
    .B1(_13009_),
    .Y(_04013_));
 sky130_fd_sc_hd__nor3b_4 _15805_ (.A(\mem_rdata_q[14] ),
    .B(\mem_rdata_q[12] ),
    .C_N(\mem_rdata_q[13] ),
    .Y(_13033_));
 sky130_fd_sc_hd__nand3_1 _15806_ (.A(_13002_),
    .B(_13019_),
    .C(_13033_),
    .Y(_13034_));
 sky130_fd_sc_hd__clkbuf_2 _15807_ (.A(_13005_),
    .X(_13035_));
 sky130_fd_sc_hd__nand2_1 _15808_ (.A(_13035_),
    .B(instr_slt),
    .Y(_13036_));
 sky130_fd_sc_hd__clkbuf_2 _15809_ (.A(_12871_),
    .X(_13037_));
 sky130_fd_sc_hd__a21oi_1 _15810_ (.A1(_13034_),
    .A2(_13036_),
    .B1(_13037_),
    .Y(_04012_));
 sky130_fd_sc_hd__nor3b_4 _15811_ (.A(_12990_),
    .B(_12991_),
    .C_N(_12993_),
    .Y(_13038_));
 sky130_fd_sc_hd__nand3_1 _15812_ (.A(_13002_),
    .B(is_alu_reg_reg),
    .C(_13038_),
    .Y(_13039_));
 sky130_fd_sc_hd__nand2_1 _15813_ (.A(_13035_),
    .B(instr_sll),
    .Y(_13040_));
 sky130_fd_sc_hd__a21oi_1 _15814_ (.A1(_13039_),
    .A2(_13040_),
    .B1(_13037_),
    .Y(_04011_));
 sky130_fd_sc_hd__nor3_4 _15815_ (.A(\mem_rdata_q[14] ),
    .B(_12991_),
    .C(_12993_),
    .Y(_13041_));
 sky130_fd_sc_hd__nand3_1 _15816_ (.A(_13018_),
    .B(is_alu_reg_reg),
    .C(_13041_),
    .Y(_13042_));
 sky130_fd_sc_hd__nand2_1 _15817_ (.A(_13035_),
    .B(instr_sub),
    .Y(_13043_));
 sky130_fd_sc_hd__a21oi_1 _15818_ (.A1(_13042_),
    .A2(_13043_),
    .B1(_13037_),
    .Y(_04010_));
 sky130_fd_sc_hd__nand3_1 _15819_ (.A(_13002_),
    .B(is_alu_reg_reg),
    .C(_13041_),
    .Y(_13044_));
 sky130_fd_sc_hd__nand2_1 _15820_ (.A(_13035_),
    .B(instr_add),
    .Y(_13045_));
 sky130_fd_sc_hd__a21oi_1 _15821_ (.A1(_13044_),
    .A2(_13045_),
    .B1(_13037_),
    .Y(_04009_));
 sky130_fd_sc_hd__clkbuf_4 _15822_ (.A(decoder_pseudo_trigger),
    .X(_13046_));
 sky130_fd_sc_hd__buf_2 _15823_ (.A(is_alu_reg_imm),
    .X(_13047_));
 sky130_fd_sc_hd__buf_4 _15824_ (.A(_12997_),
    .X(_13048_));
 sky130_fd_sc_hd__nand3b_4 _15825_ (.A_N(_13046_),
    .B(_13047_),
    .C(_13048_),
    .Y(_13049_));
 sky130_fd_sc_hd__clkbuf_4 _15826_ (.A(instr_andi),
    .X(_13050_));
 sky130_fd_sc_hd__clkbuf_2 _15827_ (.A(_13005_),
    .X(_13051_));
 sky130_fd_sc_hd__a2bb2oi_1 _15828_ (.A1_N(_12995_),
    .A2_N(_13049_),
    .B1(_13050_),
    .B2(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__nor2_1 _15829_ (.A(_12872_),
    .B(_13052_),
    .Y(_04008_));
 sky130_fd_sc_hd__buf_4 _15830_ (.A(instr_ori),
    .X(_13053_));
 sky130_fd_sc_hd__a2bb2oi_1 _15831_ (.A1_N(_13010_),
    .A2_N(_13049_),
    .B1(_13053_),
    .B2(_13051_),
    .Y(_13054_));
 sky130_fd_sc_hd__nor2_1 _15832_ (.A(_12872_),
    .B(_13054_),
    .Y(_04007_));
 sky130_vsdinv _15833_ (.A(_13049_),
    .Y(_13055_));
 sky130_fd_sc_hd__buf_2 _15834_ (.A(_13004_),
    .X(_13056_));
 sky130_fd_sc_hd__a22oi_1 _15835_ (.A1(_13055_),
    .A2(_13027_),
    .B1(instr_xori),
    .B2(_13056_),
    .Y(_13057_));
 sky130_fd_sc_hd__nor2_1 _15836_ (.A(_12872_),
    .B(_13057_),
    .Y(_04006_));
 sky130_fd_sc_hd__a22oi_1 _15837_ (.A1(_13056_),
    .A2(instr_sltiu),
    .B1(_13030_),
    .B2(_13055_),
    .Y(_13058_));
 sky130_fd_sc_hd__nor2_1 _15838_ (.A(_12872_),
    .B(_13058_),
    .Y(_04005_));
 sky130_fd_sc_hd__clkbuf_2 _15839_ (.A(_13004_),
    .X(_13059_));
 sky130_fd_sc_hd__buf_2 _15840_ (.A(_13059_),
    .X(_13060_));
 sky130_fd_sc_hd__nand2_1 _15841_ (.A(_13060_),
    .B(instr_slti),
    .Y(_13061_));
 sky130_fd_sc_hd__clkbuf_2 _15842_ (.A(_12998_),
    .X(_13062_));
 sky130_fd_sc_hd__clkbuf_2 _15843_ (.A(_13062_),
    .X(_13063_));
 sky130_fd_sc_hd__nand3_1 _15844_ (.A(_13033_),
    .B(_13047_),
    .C(_13063_),
    .Y(_13064_));
 sky130_fd_sc_hd__a21oi_1 _15845_ (.A1(_13061_),
    .A2(_13064_),
    .B1(_13037_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand2_1 _15846_ (.A(_13060_),
    .B(instr_addi),
    .Y(_13065_));
 sky130_fd_sc_hd__nand3_1 _15847_ (.A(_13041_),
    .B(_13047_),
    .C(_13063_),
    .Y(_13066_));
 sky130_fd_sc_hd__a21oi_1 _15848_ (.A1(_13065_),
    .A2(_13066_),
    .B1(_13037_),
    .Y(_04003_));
 sky130_fd_sc_hd__nand2_1 _15849_ (.A(_13051_),
    .B(instr_bgeu),
    .Y(_13067_));
 sky130_fd_sc_hd__nand3b_1 _15850_ (.A_N(_12995_),
    .B(_13063_),
    .C(_12979_),
    .Y(_13068_));
 sky130_fd_sc_hd__clkbuf_2 _15851_ (.A(_12871_),
    .X(_13069_));
 sky130_fd_sc_hd__a21oi_1 _15852_ (.A1(_13067_),
    .A2(_13068_),
    .B1(_13069_),
    .Y(_04002_));
 sky130_fd_sc_hd__clkbuf_2 _15853_ (.A(_13062_),
    .X(_13070_));
 sky130_fd_sc_hd__nand3b_1 _15854_ (.A_N(_13010_),
    .B(_12980_),
    .C(_13070_),
    .Y(_13071_));
 sky130_fd_sc_hd__nand2_1 _15855_ (.A(_13035_),
    .B(instr_bltu),
    .Y(_13072_));
 sky130_fd_sc_hd__a21oi_1 _15856_ (.A1(_13071_),
    .A2(_13072_),
    .B1(_13069_),
    .Y(_04001_));
 sky130_fd_sc_hd__nand3b_2 _15857_ (.A_N(_13020_),
    .B(_12980_),
    .C(_13070_),
    .Y(_13073_));
 sky130_fd_sc_hd__nand2_1 _15858_ (.A(_13035_),
    .B(instr_bge),
    .Y(_13074_));
 sky130_fd_sc_hd__a21oi_1 _15859_ (.A1(_13073_),
    .A2(_13074_),
    .B1(_13069_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand2_1 _15860_ (.A(_13051_),
    .B(instr_blt),
    .Y(_13075_));
 sky130_fd_sc_hd__nand3_1 _15861_ (.A(_13027_),
    .B(_12980_),
    .C(_13063_),
    .Y(_13076_));
 sky130_fd_sc_hd__a21oi_1 _15862_ (.A1(_13075_),
    .A2(_13076_),
    .B1(_13069_),
    .Y(_03999_));
 sky130_fd_sc_hd__nand2_1 _15863_ (.A(_13051_),
    .B(instr_bne),
    .Y(_13077_));
 sky130_fd_sc_hd__nand3_1 _15864_ (.A(_13038_),
    .B(_12980_),
    .C(_13063_),
    .Y(_13078_));
 sky130_fd_sc_hd__a21oi_1 _15865_ (.A1(_13077_),
    .A2(_13078_),
    .B1(_13069_),
    .Y(_03998_));
 sky130_fd_sc_hd__nand2_1 _15866_ (.A(_13051_),
    .B(instr_beq),
    .Y(_13079_));
 sky130_fd_sc_hd__nand3_1 _15867_ (.A(_13041_),
    .B(_12980_),
    .C(_13063_),
    .Y(_13080_));
 sky130_fd_sc_hd__a21oi_1 _15868_ (.A1(_13079_),
    .A2(_13080_),
    .B1(_13069_),
    .Y(_03997_));
 sky130_vsdinv _15869_ (.A(\pcpi_timeout_counter[3] ),
    .Y(_13081_));
 sky130_fd_sc_hd__nor3_4 _15870_ (.A(\pcpi_timeout_counter[2] ),
    .B(\pcpi_timeout_counter[1] ),
    .C(\pcpi_timeout_counter[0] ),
    .Y(_13082_));
 sky130_fd_sc_hd__o21ai_1 _15871_ (.A1(_13081_),
    .A2(_13082_),
    .B1(_12789_),
    .Y(_03996_));
 sky130_fd_sc_hd__o21a_1 _15872_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(\pcpi_timeout_counter[2] ),
    .X(_13083_));
 sky130_vsdinv _15873_ (.A(_12789_),
    .Y(_13084_));
 sky130_fd_sc_hd__a211o_1 _15874_ (.A1(_13082_),
    .A2(\pcpi_timeout_counter[3] ),
    .B1(_13083_),
    .C1(_13084_),
    .X(_03995_));
 sky130_fd_sc_hd__nor2_2 _15875_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .Y(_13085_));
 sky130_fd_sc_hd__o21a_1 _15876_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(\pcpi_timeout_counter[2] ),
    .B1(_13085_),
    .X(_13086_));
 sky130_fd_sc_hd__a211o_1 _15877_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(_13084_),
    .C1(_13086_),
    .X(_03994_));
 sky130_fd_sc_hd__nand3b_2 _15878_ (.A_N(\pcpi_timeout_counter[2] ),
    .B(_13085_),
    .C(_13081_),
    .Y(_13087_));
 sky130_vsdinv _15879_ (.A(_13087_),
    .Y(_13088_));
 sky130_fd_sc_hd__o21bai_1 _15880_ (.A1(\pcpi_timeout_counter[0] ),
    .A2(_13088_),
    .B1_N(_13084_),
    .Y(_03993_));
 sky130_vsdinv _15881_ (.A(mem_do_prefetch),
    .Y(_13089_));
 sky130_fd_sc_hd__a31oi_4 _15882_ (.A1(_12632_),
    .A2(net456),
    .A3(_12654_),
    .B1(_13089_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand3_1 _15883_ (.A(_12894_),
    .B(_12811_),
    .C(_12658_),
    .Y(_13090_));
 sky130_fd_sc_hd__nand3b_1 _15884_ (.A_N(_13090_),
    .B(_12920_),
    .C(_00291_),
    .Y(_13091_));
 sky130_fd_sc_hd__o2bb2ai_1 _15885_ (.A1_N(_12976_),
    .A2_N(_12890_),
    .B1(_00296_),
    .B2(_13091_),
    .Y(_03992_));
 sky130_fd_sc_hd__buf_2 _15886_ (.A(_12651_),
    .X(_13092_));
 sky130_fd_sc_hd__nand3b_2 _15887_ (.A_N(_12645_),
    .B(_12654_),
    .C(_13092_),
    .Y(_13093_));
 sky130_fd_sc_hd__o2bb2ai_1 _15888_ (.A1_N(_12645_),
    .A2_N(_12890_),
    .B1(_13093_),
    .B2(_00296_),
    .Y(_03991_));
 sky130_fd_sc_hd__buf_2 _15889_ (.A(_12848_),
    .X(_13094_));
 sky130_fd_sc_hd__clkbuf_2 _15890_ (.A(_12875_),
    .X(_13095_));
 sky130_fd_sc_hd__or2_1 _15891_ (.A(\reg_next_pc[31] ),
    .B(_13095_),
    .X(_13096_));
 sky130_fd_sc_hd__o211a_1 _15892_ (.A1(_02530_),
    .A2(_13094_),
    .B1(_12656_),
    .C1(_13096_),
    .X(_03990_));
 sky130_fd_sc_hd__buf_2 _15893_ (.A(_12876_),
    .X(_13097_));
 sky130_fd_sc_hd__or2b_1 _15894_ (.A(_02529_),
    .B_N(_12866_),
    .X(_13098_));
 sky130_fd_sc_hd__o211a_1 _15895_ (.A1(_13097_),
    .A2(\reg_next_pc[30] ),
    .B1(_12656_),
    .C1(_13098_),
    .X(_03989_));
 sky130_fd_sc_hd__clkbuf_2 _15896_ (.A(_12865_),
    .X(_13099_));
 sky130_fd_sc_hd__or2b_1 _15897_ (.A(_02527_),
    .B_N(_13099_),
    .X(_13100_));
 sky130_fd_sc_hd__o211a_1 _15898_ (.A1(_13097_),
    .A2(\reg_next_pc[29] ),
    .B1(_12656_),
    .C1(_13100_),
    .X(_03988_));
 sky130_fd_sc_hd__buf_4 _15899_ (.A(_12847_),
    .X(_13101_));
 sky130_fd_sc_hd__buf_4 _15900_ (.A(_13101_),
    .X(_00322_));
 sky130_fd_sc_hd__clkbuf_4 _15901_ (.A(_12654_),
    .X(_13102_));
 sky130_fd_sc_hd__clkbuf_2 _15902_ (.A(_13102_),
    .X(_13103_));
 sky130_vsdinv _15903_ (.A(\reg_next_pc[28] ),
    .Y(_13104_));
 sky130_fd_sc_hd__nand2_1 _15904_ (.A(_13094_),
    .B(_13104_),
    .Y(_13105_));
 sky130_fd_sc_hd__o211a_1 _15905_ (.A1(_00322_),
    .A2(_02526_),
    .B1(_13103_),
    .C1(_13105_),
    .X(_03987_));
 sky130_fd_sc_hd__or2b_1 _15906_ (.A(_02525_),
    .B_N(_13099_),
    .X(_13106_));
 sky130_fd_sc_hd__o211a_1 _15907_ (.A1(_13097_),
    .A2(\reg_next_pc[27] ),
    .B1(_13103_),
    .C1(_13106_),
    .X(_03986_));
 sky130_vsdinv _15908_ (.A(\reg_next_pc[26] ),
    .Y(_13107_));
 sky130_fd_sc_hd__nand2_1 _15909_ (.A(_13094_),
    .B(_13107_),
    .Y(_13108_));
 sky130_fd_sc_hd__o211a_1 _15910_ (.A1(_00322_),
    .A2(_02524_),
    .B1(_13103_),
    .C1(_13108_),
    .X(_03985_));
 sky130_fd_sc_hd__or2b_1 _15911_ (.A(_02523_),
    .B_N(_13099_),
    .X(_13109_));
 sky130_fd_sc_hd__o211a_1 _15912_ (.A1(_13097_),
    .A2(\reg_next_pc[25] ),
    .B1(_13103_),
    .C1(_13109_),
    .X(_03984_));
 sky130_vsdinv _15913_ (.A(\reg_next_pc[24] ),
    .Y(_13110_));
 sky130_fd_sc_hd__nand2_1 _15914_ (.A(_13094_),
    .B(_13110_),
    .Y(_13111_));
 sky130_fd_sc_hd__o211a_1 _15915_ (.A1(_00322_),
    .A2(_02522_),
    .B1(_13103_),
    .C1(_13111_),
    .X(_03983_));
 sky130_fd_sc_hd__or2b_1 _15916_ (.A(_02521_),
    .B_N(_13099_),
    .X(_13112_));
 sky130_fd_sc_hd__o211a_1 _15917_ (.A1(_13097_),
    .A2(\reg_next_pc[23] ),
    .B1(_13103_),
    .C1(_13112_),
    .X(_03982_));
 sky130_fd_sc_hd__buf_2 _15918_ (.A(_13095_),
    .X(_13113_));
 sky130_fd_sc_hd__clkbuf_2 _15919_ (.A(_13102_),
    .X(_13114_));
 sky130_fd_sc_hd__or2b_1 _15920_ (.A(_02520_),
    .B_N(_13099_),
    .X(_13115_));
 sky130_fd_sc_hd__o211a_1 _15921_ (.A1(_13113_),
    .A2(\reg_next_pc[22] ),
    .B1(_13114_),
    .C1(_13115_),
    .X(_03981_));
 sky130_fd_sc_hd__clkbuf_2 _15922_ (.A(_12848_),
    .X(_13116_));
 sky130_vsdinv _15923_ (.A(\reg_next_pc[21] ),
    .Y(_13117_));
 sky130_fd_sc_hd__nand2_1 _15924_ (.A(_13116_),
    .B(_13117_),
    .Y(_13118_));
 sky130_fd_sc_hd__o211a_1 _15925_ (.A1(_00322_),
    .A2(_02519_),
    .B1(_13114_),
    .C1(_13118_),
    .X(_03980_));
 sky130_fd_sc_hd__buf_2 _15926_ (.A(_13101_),
    .X(_13119_));
 sky130_vsdinv _15927_ (.A(\reg_next_pc[20] ),
    .Y(_13120_));
 sky130_fd_sc_hd__nand2_1 _15928_ (.A(_13116_),
    .B(_13120_),
    .Y(_13121_));
 sky130_fd_sc_hd__o211a_1 _15929_ (.A1(_13119_),
    .A2(_02518_),
    .B1(_13114_),
    .C1(_13121_),
    .X(_03979_));
 sky130_vsdinv _15930_ (.A(\reg_next_pc[19] ),
    .Y(_13122_));
 sky130_fd_sc_hd__nand2_1 _15931_ (.A(_13116_),
    .B(_13122_),
    .Y(_13123_));
 sky130_fd_sc_hd__o211a_1 _15932_ (.A1(_13119_),
    .A2(_02516_),
    .B1(_13114_),
    .C1(_13123_),
    .X(_03978_));
 sky130_fd_sc_hd__or2b_1 _15933_ (.A(_02515_),
    .B_N(_13099_),
    .X(_13124_));
 sky130_fd_sc_hd__o211a_1 _15934_ (.A1(_13113_),
    .A2(\reg_next_pc[18] ),
    .B1(_13114_),
    .C1(_13124_),
    .X(_03977_));
 sky130_vsdinv _15935_ (.A(\reg_next_pc[17] ),
    .Y(_13125_));
 sky130_fd_sc_hd__nand2_1 _15936_ (.A(_13116_),
    .B(_13125_),
    .Y(_13126_));
 sky130_fd_sc_hd__o211a_1 _15937_ (.A1(_13119_),
    .A2(_02514_),
    .B1(_13114_),
    .C1(_13126_),
    .X(_03976_));
 sky130_fd_sc_hd__buf_2 _15938_ (.A(_13102_),
    .X(_13127_));
 sky130_fd_sc_hd__clkbuf_2 _15939_ (.A(_12865_),
    .X(_13128_));
 sky130_fd_sc_hd__or2b_1 _15940_ (.A(_02513_),
    .B_N(_13128_),
    .X(_13129_));
 sky130_fd_sc_hd__o211a_1 _15941_ (.A1(_13113_),
    .A2(\reg_next_pc[16] ),
    .B1(_13127_),
    .C1(_13129_),
    .X(_03975_));
 sky130_vsdinv _15942_ (.A(\reg_next_pc[15] ),
    .Y(_13130_));
 sky130_fd_sc_hd__nand2_1 _15943_ (.A(_13116_),
    .B(_13130_),
    .Y(_13131_));
 sky130_fd_sc_hd__o211a_1 _15944_ (.A1(_13119_),
    .A2(_02512_),
    .B1(_13127_),
    .C1(_13131_),
    .X(_03974_));
 sky130_vsdinv _15945_ (.A(\reg_next_pc[14] ),
    .Y(_13132_));
 sky130_fd_sc_hd__nand2_1 _15946_ (.A(_13116_),
    .B(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__o211a_1 _15947_ (.A1(_13119_),
    .A2(_02511_),
    .B1(_13127_),
    .C1(_13133_),
    .X(_03973_));
 sky130_vsdinv _15948_ (.A(\reg_next_pc[13] ),
    .Y(_13134_));
 sky130_fd_sc_hd__nand2_1 _15949_ (.A(_12868_),
    .B(_13134_),
    .Y(_13135_));
 sky130_fd_sc_hd__o211a_1 _15950_ (.A1(_13119_),
    .A2(_02510_),
    .B1(_13127_),
    .C1(_13135_),
    .X(_03972_));
 sky130_fd_sc_hd__or2b_1 _15951_ (.A(_02509_),
    .B_N(_13128_),
    .X(_13136_));
 sky130_fd_sc_hd__o211a_1 _15952_ (.A1(_13113_),
    .A2(\reg_next_pc[12] ),
    .B1(_13127_),
    .C1(_13136_),
    .X(_03971_));
 sky130_fd_sc_hd__or2b_1 _15953_ (.A(_02508_),
    .B_N(_13128_),
    .X(_13137_));
 sky130_fd_sc_hd__o211a_1 _15954_ (.A1(_13113_),
    .A2(\reg_next_pc[11] ),
    .B1(_13127_),
    .C1(_13137_),
    .X(_03970_));
 sky130_fd_sc_hd__buf_2 _15955_ (.A(_13102_),
    .X(_13138_));
 sky130_fd_sc_hd__or2b_1 _15956_ (.A(_02507_),
    .B_N(_13128_),
    .X(_13139_));
 sky130_fd_sc_hd__o211a_1 _15957_ (.A1(_13113_),
    .A2(\reg_next_pc[10] ),
    .B1(_13138_),
    .C1(_13139_),
    .X(_03969_));
 sky130_fd_sc_hd__buf_2 _15958_ (.A(_13095_),
    .X(_13140_));
 sky130_fd_sc_hd__or2b_1 _15959_ (.A(_02537_),
    .B_N(_13128_),
    .X(_13141_));
 sky130_fd_sc_hd__o211a_1 _15960_ (.A1(_13140_),
    .A2(\reg_next_pc[9] ),
    .B1(_13138_),
    .C1(_13141_),
    .X(_03968_));
 sky130_fd_sc_hd__or2b_1 _15961_ (.A(_02536_),
    .B_N(_13128_),
    .X(_13142_));
 sky130_fd_sc_hd__o211a_1 _15962_ (.A1(_13140_),
    .A2(\reg_next_pc[8] ),
    .B1(_13138_),
    .C1(_13142_),
    .X(_03967_));
 sky130_fd_sc_hd__clkbuf_2 _15963_ (.A(_12875_),
    .X(_13143_));
 sky130_fd_sc_hd__or2b_1 _15964_ (.A(_02535_),
    .B_N(_13143_),
    .X(_13144_));
 sky130_fd_sc_hd__o211a_1 _15965_ (.A1(_13140_),
    .A2(\reg_next_pc[7] ),
    .B1(_13138_),
    .C1(_13144_),
    .X(_03966_));
 sky130_fd_sc_hd__or2b_1 _15966_ (.A(_02534_),
    .B_N(_13143_),
    .X(_13145_));
 sky130_fd_sc_hd__o211a_1 _15967_ (.A1(_13140_),
    .A2(\reg_next_pc[6] ),
    .B1(_13138_),
    .C1(_13145_),
    .X(_03965_));
 sky130_fd_sc_hd__buf_2 _15968_ (.A(_13101_),
    .X(_13146_));
 sky130_vsdinv _15969_ (.A(\reg_next_pc[5] ),
    .Y(_13147_));
 sky130_fd_sc_hd__nand2_1 _15970_ (.A(_12868_),
    .B(_13147_),
    .Y(_13148_));
 sky130_fd_sc_hd__o211a_1 _15971_ (.A1(_13146_),
    .A2(_02533_),
    .B1(_13138_),
    .C1(_13148_),
    .X(_03964_));
 sky130_fd_sc_hd__clkbuf_2 _15972_ (.A(_13102_),
    .X(_13149_));
 sky130_fd_sc_hd__or2b_1 _15973_ (.A(_02532_),
    .B_N(_13143_),
    .X(_13150_));
 sky130_fd_sc_hd__o211a_1 _15974_ (.A1(_13140_),
    .A2(\reg_next_pc[4] ),
    .B1(_13149_),
    .C1(_13150_),
    .X(_03963_));
 sky130_fd_sc_hd__or2b_1 _15975_ (.A(_02531_),
    .B_N(_13143_),
    .X(_13151_));
 sky130_fd_sc_hd__o211a_1 _15976_ (.A1(_13140_),
    .A2(\reg_next_pc[3] ),
    .B1(_13149_),
    .C1(_13151_),
    .X(_03962_));
 sky130_fd_sc_hd__clkbuf_2 _15977_ (.A(_13095_),
    .X(_13152_));
 sky130_fd_sc_hd__or2b_1 _15978_ (.A(_02528_),
    .B_N(_13143_),
    .X(_13153_));
 sky130_fd_sc_hd__o211a_1 _15979_ (.A1(_13152_),
    .A2(\reg_next_pc[2] ),
    .B1(_13149_),
    .C1(_13153_),
    .X(_03961_));
 sky130_fd_sc_hd__or2b_1 _15980_ (.A(_02517_),
    .B_N(_13143_),
    .X(_13154_));
 sky130_fd_sc_hd__o211a_1 _15981_ (.A1(_13152_),
    .A2(\reg_next_pc[1] ),
    .B1(_13149_),
    .C1(_13154_),
    .X(_03960_));
 sky130_vsdinv _15982_ (.A(\reg_pc[31] ),
    .Y(_13155_));
 sky130_fd_sc_hd__nand2_1 _15983_ (.A(_12868_),
    .B(_13155_),
    .Y(_13156_));
 sky130_fd_sc_hd__o211a_1 _15984_ (.A1(_13146_),
    .A2(_02581_),
    .B1(_13149_),
    .C1(_13156_),
    .X(_03959_));
 sky130_vsdinv _15985_ (.A(_02580_),
    .Y(_13157_));
 sky130_fd_sc_hd__nor2_1 _15986_ (.A(_12879_),
    .B(\reg_pc[30] ),
    .Y(_13158_));
 sky130_fd_sc_hd__a211oi_1 _15987_ (.A1(_13157_),
    .A2(_12877_),
    .B1(_12815_),
    .C1(_13158_),
    .Y(_03958_));
 sky130_fd_sc_hd__buf_4 _15988_ (.A(\reg_pc[29] ),
    .X(_13159_));
 sky130_fd_sc_hd__clkbuf_2 _15989_ (.A(_02579_),
    .X(_13160_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15990_ (.A(_12875_),
    .X(_13161_));
 sky130_fd_sc_hd__or2b_2 _15991_ (.A(_13160_),
    .B_N(_13161_),
    .X(_13162_));
 sky130_fd_sc_hd__o211a_1 _15992_ (.A1(_13152_),
    .A2(_13159_),
    .B1(_13149_),
    .C1(_13162_),
    .X(_03957_));
 sky130_fd_sc_hd__clkbuf_2 _15993_ (.A(_13102_),
    .X(_13163_));
 sky130_vsdinv _15994_ (.A(_02578_),
    .Y(_13164_));
 sky130_fd_sc_hd__buf_2 _15995_ (.A(_12865_),
    .X(_13165_));
 sky130_fd_sc_hd__nand2_1 _15996_ (.A(_13164_),
    .B(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__o211a_1 _15997_ (.A1(_13152_),
    .A2(\reg_pc[28] ),
    .B1(_13163_),
    .C1(_13166_),
    .X(_03956_));
 sky130_fd_sc_hd__clkbuf_2 _15998_ (.A(_02577_),
    .X(_13167_));
 sky130_vsdinv _15999_ (.A(_13167_),
    .Y(_13168_));
 sky130_fd_sc_hd__buf_6 _16000_ (.A(_12912_),
    .X(_13169_));
 sky130_fd_sc_hd__buf_4 _16001_ (.A(\reg_pc[27] ),
    .X(_13170_));
 sky130_fd_sc_hd__nor2_2 _16002_ (.A(_12879_),
    .B(_13170_),
    .Y(_13171_));
 sky130_fd_sc_hd__a211oi_4 _16003_ (.A1(_13168_),
    .A2(_12877_),
    .B1(_13169_),
    .C1(_13171_),
    .Y(_03955_));
 sky130_vsdinv _16004_ (.A(_02576_),
    .Y(_13172_));
 sky130_fd_sc_hd__buf_4 _16005_ (.A(\reg_pc[26] ),
    .X(_13173_));
 sky130_fd_sc_hd__nor2_1 _16006_ (.A(_12879_),
    .B(_13173_),
    .Y(_13174_));
 sky130_fd_sc_hd__a211oi_2 _16007_ (.A1(_13172_),
    .A2(_12877_),
    .B1(_13169_),
    .C1(_13174_),
    .Y(_03954_));
 sky130_fd_sc_hd__buf_4 _16008_ (.A(\reg_pc[25] ),
    .X(_13175_));
 sky130_fd_sc_hd__clkbuf_2 _16009_ (.A(_02575_),
    .X(_13176_));
 sky130_vsdinv _16010_ (.A(_13176_),
    .Y(_13177_));
 sky130_fd_sc_hd__nand2_1 _16011_ (.A(_13177_),
    .B(_13165_),
    .Y(_13178_));
 sky130_fd_sc_hd__o211a_1 _16012_ (.A1(_13152_),
    .A2(_13175_),
    .B1(_13163_),
    .C1(_13178_),
    .X(_03953_));
 sky130_fd_sc_hd__clkbuf_2 _16013_ (.A(_02574_),
    .X(_13179_));
 sky130_fd_sc_hd__or2b_1 _16014_ (.A(_13179_),
    .B_N(_13161_),
    .X(_13180_));
 sky130_fd_sc_hd__o211a_1 _16015_ (.A1(_13152_),
    .A2(\reg_pc[24] ),
    .B1(_13163_),
    .C1(_13180_),
    .X(_03952_));
 sky130_fd_sc_hd__clkbuf_2 _16016_ (.A(_13095_),
    .X(_13181_));
 sky130_fd_sc_hd__buf_4 _16017_ (.A(\reg_pc[23] ),
    .X(_13182_));
 sky130_fd_sc_hd__clkbuf_2 _16018_ (.A(_02573_),
    .X(_13183_));
 sky130_fd_sc_hd__or2b_1 _16019_ (.A(_13183_),
    .B_N(_13161_),
    .X(_13184_));
 sky130_fd_sc_hd__o211a_1 _16020_ (.A1(_13181_),
    .A2(_13182_),
    .B1(_13163_),
    .C1(_13184_),
    .X(_03951_));
 sky130_fd_sc_hd__buf_2 _16021_ (.A(_02572_),
    .X(_13185_));
 sky130_fd_sc_hd__clkbuf_4 _16022_ (.A(\reg_pc[22] ),
    .X(_13186_));
 sky130_fd_sc_hd__or2_1 _16023_ (.A(_12876_),
    .B(_13186_),
    .X(_13187_));
 sky130_fd_sc_hd__o211a_1 _16024_ (.A1(_13146_),
    .A2(_13185_),
    .B1(_13163_),
    .C1(_13187_),
    .X(_03950_));
 sky130_fd_sc_hd__buf_2 _16025_ (.A(_02570_),
    .X(_13188_));
 sky130_fd_sc_hd__buf_2 _16026_ (.A(\reg_pc[21] ),
    .X(_13189_));
 sky130_fd_sc_hd__or2_1 _16027_ (.A(_12876_),
    .B(_13189_),
    .X(_13190_));
 sky130_fd_sc_hd__o211a_1 _16028_ (.A1(_13146_),
    .A2(_13188_),
    .B1(_13163_),
    .C1(_13190_),
    .X(_03949_));
 sky130_vsdinv _16029_ (.A(_02569_),
    .Y(_13191_));
 sky130_fd_sc_hd__buf_2 _16030_ (.A(\reg_pc[20] ),
    .X(_13192_));
 sky130_fd_sc_hd__nor2_1 _16031_ (.A(_12866_),
    .B(_13192_),
    .Y(_13193_));
 sky130_fd_sc_hd__a211oi_1 _16032_ (.A1(_13191_),
    .A2(_12877_),
    .B1(_13169_),
    .C1(_13193_),
    .Y(_03948_));
 sky130_fd_sc_hd__buf_2 _16033_ (.A(\reg_pc[19] ),
    .X(_13194_));
 sky130_fd_sc_hd__clkbuf_4 _16034_ (.A(_12654_),
    .X(_13195_));
 sky130_fd_sc_hd__clkbuf_2 _16035_ (.A(_13195_),
    .X(_13196_));
 sky130_fd_sc_hd__clkbuf_2 _16036_ (.A(_02568_),
    .X(_13197_));
 sky130_fd_sc_hd__or2b_1 _16037_ (.A(_13197_),
    .B_N(_13161_),
    .X(_13198_));
 sky130_fd_sc_hd__o211a_1 _16038_ (.A1(_13181_),
    .A2(_13194_),
    .B1(_13196_),
    .C1(_13198_),
    .X(_03947_));
 sky130_fd_sc_hd__buf_4 _16039_ (.A(\reg_pc[18] ),
    .X(_13199_));
 sky130_fd_sc_hd__clkbuf_2 _16040_ (.A(_02567_),
    .X(_13200_));
 sky130_fd_sc_hd__or2b_1 _16041_ (.A(_13200_),
    .B_N(_13161_),
    .X(_13201_));
 sky130_fd_sc_hd__o211a_1 _16042_ (.A1(_13181_),
    .A2(_13199_),
    .B1(_13196_),
    .C1(_13201_),
    .X(_03946_));
 sky130_fd_sc_hd__clkbuf_2 _16043_ (.A(_02566_),
    .X(_13202_));
 sky130_fd_sc_hd__buf_2 _16044_ (.A(\reg_pc[17] ),
    .X(_13203_));
 sky130_fd_sc_hd__or2_1 _16045_ (.A(_12876_),
    .B(_13203_),
    .X(_13204_));
 sky130_fd_sc_hd__o211a_1 _16046_ (.A1(_13146_),
    .A2(_13202_),
    .B1(_13196_),
    .C1(_13204_),
    .X(_03945_));
 sky130_fd_sc_hd__buf_2 _16047_ (.A(\reg_pc[16] ),
    .X(_13205_));
 sky130_fd_sc_hd__clkbuf_2 _16048_ (.A(_02565_),
    .X(_13206_));
 sky130_fd_sc_hd__or2b_1 _16049_ (.A(_13206_),
    .B_N(_13161_),
    .X(_13207_));
 sky130_fd_sc_hd__o211a_1 _16050_ (.A1(_13181_),
    .A2(_13205_),
    .B1(_13196_),
    .C1(_13207_),
    .X(_03944_));
 sky130_fd_sc_hd__buf_2 _16051_ (.A(\reg_pc[15] ),
    .X(_13208_));
 sky130_fd_sc_hd__clkbuf_2 _16052_ (.A(_02564_),
    .X(_13209_));
 sky130_fd_sc_hd__clkbuf_2 _16053_ (.A(_12875_),
    .X(_13210_));
 sky130_fd_sc_hd__or2b_1 _16054_ (.A(_13209_),
    .B_N(_13210_),
    .X(_13211_));
 sky130_fd_sc_hd__o211a_1 _16055_ (.A1(_13181_),
    .A2(_13208_),
    .B1(_13196_),
    .C1(_13211_),
    .X(_03943_));
 sky130_vsdinv _16056_ (.A(_02563_),
    .Y(_13212_));
 sky130_fd_sc_hd__buf_2 _16057_ (.A(\reg_pc[14] ),
    .X(_13213_));
 sky130_fd_sc_hd__nor2_1 _16058_ (.A(_12866_),
    .B(_13213_),
    .Y(_13214_));
 sky130_fd_sc_hd__a211oi_2 _16059_ (.A1(_13212_),
    .A2(_13097_),
    .B1(_13169_),
    .C1(_13214_),
    .Y(_03942_));
 sky130_fd_sc_hd__buf_2 _16060_ (.A(\reg_pc[13] ),
    .X(_13215_));
 sky130_fd_sc_hd__clkbuf_2 _16061_ (.A(_02562_),
    .X(_13216_));
 sky130_fd_sc_hd__or2b_1 _16062_ (.A(_13216_),
    .B_N(_13210_),
    .X(_13217_));
 sky130_fd_sc_hd__o211a_1 _16063_ (.A1(_13181_),
    .A2(_13215_),
    .B1(_13196_),
    .C1(_13217_),
    .X(_03941_));
 sky130_fd_sc_hd__clkbuf_2 _16064_ (.A(_02561_),
    .X(_13218_));
 sky130_fd_sc_hd__clkbuf_2 _16065_ (.A(_13195_),
    .X(_13219_));
 sky130_fd_sc_hd__inv_2 _16066_ (.A(\reg_pc[12] ),
    .Y(_13220_));
 sky130_fd_sc_hd__nand2_1 _16067_ (.A(_12868_),
    .B(_13220_),
    .Y(_13221_));
 sky130_fd_sc_hd__o211a_1 _16068_ (.A1(_13146_),
    .A2(_13218_),
    .B1(_13219_),
    .C1(_13221_),
    .X(_03940_));
 sky130_fd_sc_hd__clkbuf_2 _16069_ (.A(_12865_),
    .X(_13222_));
 sky130_fd_sc_hd__clkbuf_4 _16070_ (.A(\reg_pc[11] ),
    .X(_13223_));
 sky130_fd_sc_hd__clkbuf_2 _16071_ (.A(_02589_),
    .X(_13224_));
 sky130_fd_sc_hd__or2b_1 _16072_ (.A(_13224_),
    .B_N(_13210_),
    .X(_13225_));
 sky130_fd_sc_hd__o211a_1 _16073_ (.A1(_13222_),
    .A2(_13223_),
    .B1(_13219_),
    .C1(_13225_),
    .X(_03939_));
 sky130_fd_sc_hd__buf_2 _16074_ (.A(\reg_pc[10] ),
    .X(_13226_));
 sky130_fd_sc_hd__clkbuf_2 _16075_ (.A(_02588_),
    .X(_13227_));
 sky130_fd_sc_hd__or2b_1 _16076_ (.A(_13227_),
    .B_N(_13210_),
    .X(_13228_));
 sky130_fd_sc_hd__o211a_1 _16077_ (.A1(_13222_),
    .A2(_13226_),
    .B1(_13219_),
    .C1(_13228_),
    .X(_03938_));
 sky130_fd_sc_hd__clkbuf_2 _16078_ (.A(\reg_pc[9] ),
    .X(_13229_));
 sky130_fd_sc_hd__clkbuf_2 _16079_ (.A(_02587_),
    .X(_13230_));
 sky130_fd_sc_hd__or2b_1 _16080_ (.A(_13230_),
    .B_N(_13210_),
    .X(_13231_));
 sky130_fd_sc_hd__o211a_1 _16081_ (.A1(_13222_),
    .A2(_13229_),
    .B1(_13219_),
    .C1(_13231_),
    .X(_03937_));
 sky130_fd_sc_hd__clkbuf_2 _16082_ (.A(_02586_),
    .X(_13232_));
 sky130_fd_sc_hd__inv_2 _16083_ (.A(\reg_pc[8] ),
    .Y(_13233_));
 sky130_fd_sc_hd__nand2_1 _16084_ (.A(_12868_),
    .B(_13233_),
    .Y(_13234_));
 sky130_fd_sc_hd__o211a_1 _16085_ (.A1(_13094_),
    .A2(_13232_),
    .B1(_13219_),
    .C1(_13234_),
    .X(_03936_));
 sky130_vsdinv _16086_ (.A(_02585_),
    .Y(_13235_));
 sky130_fd_sc_hd__nand2_1 _16087_ (.A(_13235_),
    .B(_13165_),
    .Y(_13236_));
 sky130_fd_sc_hd__o211a_1 _16088_ (.A1(_13222_),
    .A2(\reg_pc[7] ),
    .B1(_13219_),
    .C1(_13236_),
    .X(_03935_));
 sky130_fd_sc_hd__clkbuf_4 _16089_ (.A(\reg_pc[6] ),
    .X(_13237_));
 sky130_fd_sc_hd__buf_4 _16090_ (.A(_13195_),
    .X(_13238_));
 sky130_fd_sc_hd__clkbuf_2 _16091_ (.A(_02584_),
    .X(_13239_));
 sky130_fd_sc_hd__or2b_1 _16092_ (.A(_13239_),
    .B_N(_13210_),
    .X(_13240_));
 sky130_fd_sc_hd__o211a_1 _16093_ (.A1(_13222_),
    .A2(_13237_),
    .B1(_13238_),
    .C1(_13240_),
    .X(_03934_));
 sky130_fd_sc_hd__clkbuf_4 _16094_ (.A(\reg_pc[5] ),
    .X(_13241_));
 sky130_vsdinv _16095_ (.A(_02583_),
    .Y(_13242_));
 sky130_fd_sc_hd__nand2_1 _16096_ (.A(_13242_),
    .B(_13165_),
    .Y(_13243_));
 sky130_fd_sc_hd__o211a_1 _16097_ (.A1(_13222_),
    .A2(_13241_),
    .B1(_13238_),
    .C1(_13243_),
    .X(_03933_));
 sky130_fd_sc_hd__clkbuf_4 _16098_ (.A(\reg_pc[4] ),
    .X(_13244_));
 sky130_fd_sc_hd__nor2_1 _16099_ (.A(_12866_),
    .B(_13244_),
    .Y(_13245_));
 sky130_fd_sc_hd__a211oi_2 _16100_ (.A1(_12877_),
    .A2(_01475_),
    .B1(_13169_),
    .C1(_13245_),
    .Y(_03932_));
 sky130_fd_sc_hd__inv_2 _16101_ (.A(_01475_),
    .Y(_02582_));
 sky130_fd_sc_hd__buf_2 _16102_ (.A(\reg_pc[3] ),
    .X(_13246_));
 sky130_fd_sc_hd__clkbuf_2 _16103_ (.A(_02571_),
    .X(_13247_));
 sky130_fd_sc_hd__or2b_1 _16104_ (.A(_13247_),
    .B_N(_12876_),
    .X(_13248_));
 sky130_fd_sc_hd__o211a_1 _16105_ (.A1(_13165_),
    .A2(_13246_),
    .B1(_13238_),
    .C1(_13248_),
    .X(_03931_));
 sky130_fd_sc_hd__buf_2 _16106_ (.A(\reg_pc[2] ),
    .X(_13249_));
 sky130_fd_sc_hd__buf_2 _16107_ (.A(_02560_),
    .X(_13250_));
 sky130_fd_sc_hd__inv_2 _16108_ (.A(_13250_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_1 _16109_ (.A(_01561_),
    .B(_12879_),
    .Y(_13251_));
 sky130_fd_sc_hd__o211a_1 _16110_ (.A1(_13165_),
    .A2(_13249_),
    .B1(_13238_),
    .C1(_13251_),
    .X(_03930_));
 sky130_fd_sc_hd__or2_1 _16111_ (.A(_13095_),
    .B(\reg_pc[1] ),
    .X(_13252_));
 sky130_fd_sc_hd__o211a_1 _16112_ (.A1(_13094_),
    .A2(_02590_),
    .B1(_13238_),
    .C1(_13252_),
    .X(_03929_));
 sky130_vsdinv _16113_ (.A(\count_instr[63] ),
    .Y(_13253_));
 sky130_vsdinv _16114_ (.A(\count_instr[58] ),
    .Y(_13254_));
 sky130_vsdinv _16115_ (.A(\count_instr[57] ),
    .Y(_13255_));
 sky130_vsdinv _16116_ (.A(\count_instr[54] ),
    .Y(_13256_));
 sky130_vsdinv _16117_ (.A(\count_instr[53] ),
    .Y(_13257_));
 sky130_vsdinv _16118_ (.A(\count_instr[50] ),
    .Y(_13258_));
 sky130_vsdinv _16119_ (.A(\count_instr[49] ),
    .Y(_13259_));
 sky130_vsdinv _16120_ (.A(\count_instr[46] ),
    .Y(_13260_));
 sky130_vsdinv _16121_ (.A(\count_instr[45] ),
    .Y(_13261_));
 sky130_vsdinv _16122_ (.A(\count_instr[42] ),
    .Y(_13262_));
 sky130_vsdinv _16123_ (.A(\count_instr[41] ),
    .Y(_13263_));
 sky130_vsdinv _16124_ (.A(\count_instr[38] ),
    .Y(_13264_));
 sky130_vsdinv _16125_ (.A(\count_instr[37] ),
    .Y(_13265_));
 sky130_fd_sc_hd__inv_2 _16126_ (.A(\count_instr[34] ),
    .Y(_13266_));
 sky130_fd_sc_hd__inv_2 _16127_ (.A(\count_instr[33] ),
    .Y(_13267_));
 sky130_vsdinv _16128_ (.A(\count_instr[30] ),
    .Y(_13268_));
 sky130_vsdinv _16129_ (.A(\count_instr[29] ),
    .Y(_13269_));
 sky130_fd_sc_hd__inv_2 _16130_ (.A(\count_instr[26] ),
    .Y(_13270_));
 sky130_fd_sc_hd__inv_2 _16131_ (.A(\count_instr[25] ),
    .Y(_13271_));
 sky130_fd_sc_hd__inv_2 _16132_ (.A(\count_instr[22] ),
    .Y(_13272_));
 sky130_fd_sc_hd__inv_2 _16133_ (.A(\count_instr[21] ),
    .Y(_13273_));
 sky130_fd_sc_hd__inv_2 _16134_ (.A(\count_instr[18] ),
    .Y(_13274_));
 sky130_fd_sc_hd__inv_2 _16135_ (.A(\count_instr[17] ),
    .Y(_13275_));
 sky130_vsdinv _16136_ (.A(\count_instr[14] ),
    .Y(_13276_));
 sky130_vsdinv _16137_ (.A(\count_instr[13] ),
    .Y(_13277_));
 sky130_vsdinv _16138_ (.A(\count_instr[10] ),
    .Y(_13278_));
 sky130_vsdinv _16139_ (.A(\count_instr[9] ),
    .Y(_13279_));
 sky130_fd_sc_hd__inv_2 _16140_ (.A(\count_instr[6] ),
    .Y(_13280_));
 sky130_fd_sc_hd__inv_2 _16141_ (.A(\count_instr[5] ),
    .Y(_13281_));
 sky130_vsdinv _16142_ (.A(\count_instr[0] ),
    .Y(_13282_));
 sky130_fd_sc_hd__and2_1 _16143_ (.A(\count_instr[2] ),
    .B(\count_instr[1] ),
    .X(_13283_));
 sky130_vsdinv _16144_ (.A(_13283_),
    .Y(_13284_));
 sky130_fd_sc_hd__nor3_4 _16145_ (.A(_13282_),
    .B(_13284_),
    .C(_12772_),
    .Y(_13285_));
 sky130_fd_sc_hd__nand3_4 _16146_ (.A(_13285_),
    .B(\count_instr[4] ),
    .C(\count_instr[3] ),
    .Y(_13286_));
 sky130_fd_sc_hd__nor3_4 _16147_ (.A(_13280_),
    .B(_13281_),
    .C(_13286_),
    .Y(_13287_));
 sky130_fd_sc_hd__nand3_4 _16148_ (.A(_13287_),
    .B(\count_instr[8] ),
    .C(\count_instr[7] ),
    .Y(_13288_));
 sky130_fd_sc_hd__nor3_4 _16149_ (.A(_13278_),
    .B(_13279_),
    .C(_13288_),
    .Y(_13289_));
 sky130_fd_sc_hd__nand3_4 _16150_ (.A(_13289_),
    .B(\count_instr[12] ),
    .C(\count_instr[11] ),
    .Y(_13290_));
 sky130_fd_sc_hd__nor3_4 _16151_ (.A(_13276_),
    .B(_13277_),
    .C(_13290_),
    .Y(_13291_));
 sky130_fd_sc_hd__nand3_4 _16152_ (.A(_13291_),
    .B(\count_instr[16] ),
    .C(\count_instr[15] ),
    .Y(_13292_));
 sky130_fd_sc_hd__nor3_4 _16153_ (.A(_13274_),
    .B(_13275_),
    .C(_13292_),
    .Y(_13293_));
 sky130_fd_sc_hd__nand3_4 _16154_ (.A(_13293_),
    .B(\count_instr[20] ),
    .C(\count_instr[19] ),
    .Y(_13294_));
 sky130_fd_sc_hd__nor3_4 _16155_ (.A(_13272_),
    .B(_13273_),
    .C(_13294_),
    .Y(_13295_));
 sky130_fd_sc_hd__nand3_4 _16156_ (.A(_13295_),
    .B(\count_instr[24] ),
    .C(\count_instr[23] ),
    .Y(_13296_));
 sky130_fd_sc_hd__nor3_4 _16157_ (.A(_13270_),
    .B(_13271_),
    .C(_13296_),
    .Y(_13297_));
 sky130_fd_sc_hd__nand3_4 _16158_ (.A(_13297_),
    .B(\count_instr[28] ),
    .C(\count_instr[27] ),
    .Y(_13298_));
 sky130_fd_sc_hd__nor3_4 _16159_ (.A(_13268_),
    .B(_13269_),
    .C(_13298_),
    .Y(_13299_));
 sky130_fd_sc_hd__nand3_4 _16160_ (.A(_13299_),
    .B(\count_instr[32] ),
    .C(\count_instr[31] ),
    .Y(_13300_));
 sky130_fd_sc_hd__nor3_4 _16161_ (.A(_13266_),
    .B(_13267_),
    .C(_13300_),
    .Y(_13301_));
 sky130_fd_sc_hd__nand3_4 _16162_ (.A(_13301_),
    .B(\count_instr[36] ),
    .C(\count_instr[35] ),
    .Y(_13302_));
 sky130_fd_sc_hd__nor3_4 _16163_ (.A(_13264_),
    .B(_13265_),
    .C(_13302_),
    .Y(_13303_));
 sky130_fd_sc_hd__nand3_4 _16164_ (.A(_13303_),
    .B(\count_instr[40] ),
    .C(\count_instr[39] ),
    .Y(_13304_));
 sky130_fd_sc_hd__nor3_4 _16165_ (.A(_13262_),
    .B(_13263_),
    .C(_13304_),
    .Y(_13305_));
 sky130_fd_sc_hd__nand3_4 _16166_ (.A(_13305_),
    .B(\count_instr[44] ),
    .C(\count_instr[43] ),
    .Y(_13306_));
 sky130_fd_sc_hd__nor3_4 _16167_ (.A(_13260_),
    .B(_13261_),
    .C(_13306_),
    .Y(_13307_));
 sky130_fd_sc_hd__nand3_4 _16168_ (.A(_13307_),
    .B(\count_instr[48] ),
    .C(\count_instr[47] ),
    .Y(_13308_));
 sky130_fd_sc_hd__nor3_4 _16169_ (.A(_13258_),
    .B(_13259_),
    .C(_13308_),
    .Y(_13309_));
 sky130_fd_sc_hd__nand3_4 _16170_ (.A(_13309_),
    .B(\count_instr[52] ),
    .C(\count_instr[51] ),
    .Y(_13310_));
 sky130_fd_sc_hd__nor3_4 _16171_ (.A(_13256_),
    .B(_13257_),
    .C(_13310_),
    .Y(_13311_));
 sky130_fd_sc_hd__nand3_4 _16172_ (.A(_13311_),
    .B(\count_instr[56] ),
    .C(\count_instr[55] ),
    .Y(_13312_));
 sky130_fd_sc_hd__nor3_4 _16173_ (.A(_13254_),
    .B(_13255_),
    .C(_13312_),
    .Y(_13313_));
 sky130_fd_sc_hd__nand3_4 _16174_ (.A(_13313_),
    .B(\count_instr[60] ),
    .C(\count_instr[59] ),
    .Y(_13314_));
 sky130_fd_sc_hd__nand3b_1 _16175_ (.A_N(_13314_),
    .B(\count_instr[62] ),
    .C(\count_instr[61] ),
    .Y(_13315_));
 sky130_fd_sc_hd__nor2_1 _16176_ (.A(_13253_),
    .B(_13315_),
    .Y(_13316_));
 sky130_vsdinv _16177_ (.A(\count_instr[62] ),
    .Y(_13317_));
 sky130_vsdinv _16178_ (.A(\count_instr[61] ),
    .Y(_13318_));
 sky130_fd_sc_hd__nor3_4 _16179_ (.A(_13317_),
    .B(_13318_),
    .C(_13314_),
    .Y(_13319_));
 sky130_fd_sc_hd__o21bai_1 _16180_ (.A1(\count_instr[63] ),
    .A2(_13319_),
    .B1_N(_12814_),
    .Y(_13320_));
 sky130_fd_sc_hd__nor2_1 _16181_ (.A(_13316_),
    .B(_13320_),
    .Y(_03928_));
 sky130_fd_sc_hd__clkbuf_2 _16182_ (.A(_12643_),
    .X(_13321_));
 sky130_fd_sc_hd__buf_4 _16183_ (.A(_13321_),
    .X(_13322_));
 sky130_fd_sc_hd__a41oi_1 _16184_ (.A1(\count_instr[61] ),
    .A2(_13313_),
    .A3(\count_instr[60] ),
    .A4(\count_instr[59] ),
    .B1(\count_instr[62] ),
    .Y(_13323_));
 sky130_fd_sc_hd__nor3_1 _16185_ (.A(_13322_),
    .B(_13323_),
    .C(_13319_),
    .Y(_03927_));
 sky130_fd_sc_hd__o21bai_1 _16186_ (.A1(_13318_),
    .A2(_13314_),
    .B1_N(_12814_),
    .Y(_13324_));
 sky130_fd_sc_hd__a21oi_1 _16187_ (.A1(_13318_),
    .A2(_13314_),
    .B1(_13324_),
    .Y(_03926_));
 sky130_vsdinv _16188_ (.A(\count_instr[59] ),
    .Y(_13325_));
 sky130_fd_sc_hd__nand3b_2 _16189_ (.A_N(_13312_),
    .B(\count_instr[58] ),
    .C(\count_instr[57] ),
    .Y(_13326_));
 sky130_fd_sc_hd__nor2_1 _16190_ (.A(_13325_),
    .B(_13326_),
    .Y(_13327_));
 sky130_fd_sc_hd__a31oi_1 _16191_ (.A1(_13313_),
    .A2(\count_instr[60] ),
    .A3(\count_instr[59] ),
    .B1(_12964_),
    .Y(_13328_));
 sky130_fd_sc_hd__o21a_1 _16192_ (.A1(\count_instr[60] ),
    .A2(_13327_),
    .B1(_13328_),
    .X(_03925_));
 sky130_fd_sc_hd__clkbuf_4 _16193_ (.A(_12895_),
    .X(_13329_));
 sky130_fd_sc_hd__o41ai_1 _16194_ (.A1(_13325_),
    .A2(_13254_),
    .A3(_13255_),
    .A4(_13312_),
    .B1(_13329_),
    .Y(_13330_));
 sky130_fd_sc_hd__a21oi_1 _16195_ (.A1(_13325_),
    .A2(_13326_),
    .B1(_13330_),
    .Y(_03924_));
 sky130_fd_sc_hd__nor2_1 _16196_ (.A(_13255_),
    .B(_13312_),
    .Y(_13331_));
 sky130_vsdinv _16197_ (.A(_13331_),
    .Y(_13332_));
 sky130_fd_sc_hd__buf_4 _16198_ (.A(_12895_),
    .X(_13333_));
 sky130_fd_sc_hd__o31ai_1 _16199_ (.A1(_13254_),
    .A2(_13255_),
    .A3(_13312_),
    .B1(_13333_),
    .Y(_13334_));
 sky130_fd_sc_hd__a21oi_1 _16200_ (.A1(_13332_),
    .A2(_13254_),
    .B1(_13334_),
    .Y(_03923_));
 sky130_fd_sc_hd__a31oi_1 _16201_ (.A1(_13311_),
    .A2(\count_instr[56] ),
    .A3(\count_instr[55] ),
    .B1(\count_instr[57] ),
    .Y(_13335_));
 sky130_fd_sc_hd__nor3_1 _16202_ (.A(_13322_),
    .B(_13335_),
    .C(_13331_),
    .Y(_03922_));
 sky130_vsdinv _16203_ (.A(\count_instr[55] ),
    .Y(_13336_));
 sky130_vsdinv _16204_ (.A(\count_instr[51] ),
    .Y(_13337_));
 sky130_vsdinv _16205_ (.A(\count_instr[47] ),
    .Y(_13338_));
 sky130_vsdinv _16206_ (.A(\count_instr[43] ),
    .Y(_13339_));
 sky130_vsdinv _16207_ (.A(\count_instr[39] ),
    .Y(_13340_));
 sky130_vsdinv _16208_ (.A(\count_instr[35] ),
    .Y(_13341_));
 sky130_vsdinv _16209_ (.A(\count_instr[31] ),
    .Y(_13342_));
 sky130_vsdinv _16210_ (.A(\count_instr[27] ),
    .Y(_13343_));
 sky130_vsdinv _16211_ (.A(\count_instr[23] ),
    .Y(_13344_));
 sky130_vsdinv _16212_ (.A(\count_instr[19] ),
    .Y(_13345_));
 sky130_vsdinv _16213_ (.A(\count_instr[15] ),
    .Y(_13346_));
 sky130_vsdinv _16214_ (.A(\count_instr[11] ),
    .Y(_13347_));
 sky130_vsdinv _16215_ (.A(\count_instr[7] ),
    .Y(_13348_));
 sky130_fd_sc_hd__and4_1 _16216_ (.A(_12773_),
    .B(\count_instr[3] ),
    .C(\count_instr[0] ),
    .D(_13283_),
    .X(_13349_));
 sky130_fd_sc_hd__nand3_4 _16217_ (.A(_13349_),
    .B(\count_instr[5] ),
    .C(\count_instr[4] ),
    .Y(_13350_));
 sky130_fd_sc_hd__nor3_4 _16218_ (.A(_13348_),
    .B(_13280_),
    .C(_13350_),
    .Y(_13351_));
 sky130_fd_sc_hd__nand3_2 _16219_ (.A(_13351_),
    .B(\count_instr[9] ),
    .C(\count_instr[8] ),
    .Y(_13352_));
 sky130_fd_sc_hd__nor3_4 _16220_ (.A(_13347_),
    .B(_13278_),
    .C(_13352_),
    .Y(_13353_));
 sky130_fd_sc_hd__nand3_2 _16221_ (.A(_13353_),
    .B(\count_instr[13] ),
    .C(\count_instr[12] ),
    .Y(_13354_));
 sky130_fd_sc_hd__nor3_4 _16222_ (.A(_13346_),
    .B(_13276_),
    .C(_13354_),
    .Y(_13355_));
 sky130_fd_sc_hd__nand3_4 _16223_ (.A(_13355_),
    .B(\count_instr[17] ),
    .C(\count_instr[16] ),
    .Y(_13356_));
 sky130_fd_sc_hd__nor3_4 _16224_ (.A(_13345_),
    .B(_13274_),
    .C(_13356_),
    .Y(_13357_));
 sky130_fd_sc_hd__nand3_4 _16225_ (.A(_13357_),
    .B(\count_instr[21] ),
    .C(\count_instr[20] ),
    .Y(_13358_));
 sky130_fd_sc_hd__nor3_4 _16226_ (.A(_13344_),
    .B(_13272_),
    .C(_13358_),
    .Y(_13359_));
 sky130_fd_sc_hd__nand3_4 _16227_ (.A(_13359_),
    .B(\count_instr[25] ),
    .C(\count_instr[24] ),
    .Y(_13360_));
 sky130_fd_sc_hd__nor3_4 _16228_ (.A(_13343_),
    .B(_13270_),
    .C(_13360_),
    .Y(_13361_));
 sky130_fd_sc_hd__nand3_2 _16229_ (.A(_13361_),
    .B(\count_instr[29] ),
    .C(\count_instr[28] ),
    .Y(_13362_));
 sky130_fd_sc_hd__nor3_4 _16230_ (.A(_13342_),
    .B(_13268_),
    .C(_13362_),
    .Y(_13363_));
 sky130_fd_sc_hd__nand3_4 _16231_ (.A(_13363_),
    .B(\count_instr[33] ),
    .C(\count_instr[32] ),
    .Y(_13364_));
 sky130_fd_sc_hd__nor3_4 _16232_ (.A(_13341_),
    .B(_13266_),
    .C(_13364_),
    .Y(_13365_));
 sky130_fd_sc_hd__nand3_2 _16233_ (.A(_13365_),
    .B(\count_instr[37] ),
    .C(\count_instr[36] ),
    .Y(_13366_));
 sky130_fd_sc_hd__nor3_4 _16234_ (.A(_13340_),
    .B(_13264_),
    .C(_13366_),
    .Y(_13367_));
 sky130_fd_sc_hd__nand3_2 _16235_ (.A(_13367_),
    .B(\count_instr[41] ),
    .C(\count_instr[40] ),
    .Y(_13368_));
 sky130_fd_sc_hd__nor3_4 _16236_ (.A(_13339_),
    .B(_13262_),
    .C(_13368_),
    .Y(_13369_));
 sky130_fd_sc_hd__nand3_2 _16237_ (.A(_13369_),
    .B(\count_instr[45] ),
    .C(\count_instr[44] ),
    .Y(_13370_));
 sky130_fd_sc_hd__nor3_4 _16238_ (.A(_13338_),
    .B(_13260_),
    .C(_13370_),
    .Y(_13371_));
 sky130_fd_sc_hd__nand3_2 _16239_ (.A(_13371_),
    .B(\count_instr[49] ),
    .C(\count_instr[48] ),
    .Y(_13372_));
 sky130_fd_sc_hd__nor3_4 _16240_ (.A(_13337_),
    .B(_13258_),
    .C(_13372_),
    .Y(_13373_));
 sky130_fd_sc_hd__nand3_2 _16241_ (.A(_13373_),
    .B(\count_instr[53] ),
    .C(\count_instr[52] ),
    .Y(_13374_));
 sky130_fd_sc_hd__nor3_2 _16242_ (.A(_13336_),
    .B(_13256_),
    .C(_13374_),
    .Y(_13375_));
 sky130_fd_sc_hd__a31oi_1 _16243_ (.A1(_13311_),
    .A2(\count_instr[56] ),
    .A3(\count_instr[55] ),
    .B1(_12964_),
    .Y(_13376_));
 sky130_fd_sc_hd__o21a_1 _16244_ (.A1(\count_instr[56] ),
    .A2(_13375_),
    .B1(_13376_),
    .X(_03921_));
 sky130_vsdinv _16245_ (.A(_13311_),
    .Y(_13377_));
 sky130_fd_sc_hd__o41ai_1 _16246_ (.A1(_13336_),
    .A2(_13256_),
    .A3(_13257_),
    .A4(_13310_),
    .B1(_13329_),
    .Y(_13378_));
 sky130_fd_sc_hd__a21oi_1 _16247_ (.A1(_13336_),
    .A2(_13377_),
    .B1(_13378_),
    .Y(_03920_));
 sky130_fd_sc_hd__a41oi_1 _16248_ (.A1(\count_instr[53] ),
    .A2(_13309_),
    .A3(\count_instr[52] ),
    .A4(\count_instr[51] ),
    .B1(\count_instr[54] ),
    .Y(_13379_));
 sky130_fd_sc_hd__nor3_1 _16249_ (.A(_13322_),
    .B(_13379_),
    .C(_13311_),
    .Y(_03919_));
 sky130_fd_sc_hd__o21bai_1 _16250_ (.A1(_13257_),
    .A2(_13310_),
    .B1_N(_12814_),
    .Y(_13380_));
 sky130_fd_sc_hd__a21oi_1 _16251_ (.A1(_13257_),
    .A2(_13310_),
    .B1(_13380_),
    .Y(_03918_));
 sky130_fd_sc_hd__a31oi_1 _16252_ (.A1(_13309_),
    .A2(\count_instr[52] ),
    .A3(\count_instr[51] ),
    .B1(_12964_),
    .Y(_13381_));
 sky130_fd_sc_hd__o21a_1 _16253_ (.A1(\count_instr[52] ),
    .A2(_13373_),
    .B1(_13381_),
    .X(_03917_));
 sky130_vsdinv _16254_ (.A(_13309_),
    .Y(_13382_));
 sky130_fd_sc_hd__buf_2 _16255_ (.A(_12895_),
    .X(_13383_));
 sky130_fd_sc_hd__o41ai_1 _16256_ (.A1(_13337_),
    .A2(_13258_),
    .A3(_13259_),
    .A4(_13308_),
    .B1(_13383_),
    .Y(_13384_));
 sky130_fd_sc_hd__a21oi_1 _16257_ (.A1(_13337_),
    .A2(_13382_),
    .B1(_13384_),
    .Y(_03916_));
 sky130_fd_sc_hd__a41oi_1 _16258_ (.A1(\count_instr[49] ),
    .A2(_13307_),
    .A3(\count_instr[48] ),
    .A4(\count_instr[47] ),
    .B1(\count_instr[50] ),
    .Y(_13385_));
 sky130_fd_sc_hd__nor3_1 _16259_ (.A(_13322_),
    .B(_13385_),
    .C(_13309_),
    .Y(_03915_));
 sky130_fd_sc_hd__clkbuf_2 _16260_ (.A(_12643_),
    .X(_13386_));
 sky130_fd_sc_hd__o21bai_1 _16261_ (.A1(_13259_),
    .A2(_13308_),
    .B1_N(_13386_),
    .Y(_13387_));
 sky130_fd_sc_hd__a21oi_1 _16262_ (.A1(_13259_),
    .A2(_13308_),
    .B1(_13387_),
    .Y(_03914_));
 sky130_fd_sc_hd__buf_2 _16263_ (.A(_12912_),
    .X(_13388_));
 sky130_fd_sc_hd__a31oi_1 _16264_ (.A1(_13307_),
    .A2(\count_instr[48] ),
    .A3(\count_instr[47] ),
    .B1(_13388_),
    .Y(_13389_));
 sky130_fd_sc_hd__o21a_1 _16265_ (.A1(\count_instr[48] ),
    .A2(_13371_),
    .B1(_13389_),
    .X(_03913_));
 sky130_vsdinv _16266_ (.A(_13307_),
    .Y(_13390_));
 sky130_fd_sc_hd__o41ai_1 _16267_ (.A1(_13338_),
    .A2(_13260_),
    .A3(_13261_),
    .A4(_13306_),
    .B1(_13383_),
    .Y(_13391_));
 sky130_fd_sc_hd__a21oi_1 _16268_ (.A1(_13338_),
    .A2(_13390_),
    .B1(_13391_),
    .Y(_03912_));
 sky130_fd_sc_hd__buf_2 _16269_ (.A(_13321_),
    .X(_13392_));
 sky130_fd_sc_hd__a41oi_1 _16270_ (.A1(\count_instr[45] ),
    .A2(_13305_),
    .A3(\count_instr[44] ),
    .A4(\count_instr[43] ),
    .B1(\count_instr[46] ),
    .Y(_13393_));
 sky130_fd_sc_hd__nor3_1 _16271_ (.A(_13392_),
    .B(_13393_),
    .C(_13307_),
    .Y(_03911_));
 sky130_fd_sc_hd__o21bai_1 _16272_ (.A1(_13261_),
    .A2(_13306_),
    .B1_N(_13386_),
    .Y(_13394_));
 sky130_fd_sc_hd__a21oi_1 _16273_ (.A1(_13261_),
    .A2(_13306_),
    .B1(_13394_),
    .Y(_03910_));
 sky130_fd_sc_hd__a31oi_1 _16274_ (.A1(_13305_),
    .A2(\count_instr[44] ),
    .A3(\count_instr[43] ),
    .B1(_13388_),
    .Y(_13395_));
 sky130_fd_sc_hd__o21a_1 _16275_ (.A1(\count_instr[44] ),
    .A2(_13369_),
    .B1(_13395_),
    .X(_03909_));
 sky130_vsdinv _16276_ (.A(_13305_),
    .Y(_13396_));
 sky130_fd_sc_hd__o41ai_1 _16277_ (.A1(_13339_),
    .A2(_13262_),
    .A3(_13263_),
    .A4(_13304_),
    .B1(_13383_),
    .Y(_13397_));
 sky130_fd_sc_hd__a21oi_1 _16278_ (.A1(_13339_),
    .A2(_13396_),
    .B1(_13397_),
    .Y(_03908_));
 sky130_fd_sc_hd__a41oi_1 _16279_ (.A1(\count_instr[41] ),
    .A2(_13303_),
    .A3(\count_instr[40] ),
    .A4(\count_instr[39] ),
    .B1(\count_instr[42] ),
    .Y(_13398_));
 sky130_fd_sc_hd__nor3_1 _16280_ (.A(_13392_),
    .B(_13398_),
    .C(_13305_),
    .Y(_03907_));
 sky130_fd_sc_hd__o21bai_1 _16281_ (.A1(_13263_),
    .A2(_13304_),
    .B1_N(_13386_),
    .Y(_13399_));
 sky130_fd_sc_hd__a21oi_1 _16282_ (.A1(_13263_),
    .A2(_13304_),
    .B1(_13399_),
    .Y(_03906_));
 sky130_fd_sc_hd__a31oi_1 _16283_ (.A1(_13303_),
    .A2(\count_instr[40] ),
    .A3(\count_instr[39] ),
    .B1(_13388_),
    .Y(_13400_));
 sky130_fd_sc_hd__o21a_1 _16284_ (.A1(\count_instr[40] ),
    .A2(_13367_),
    .B1(_13400_),
    .X(_03905_));
 sky130_vsdinv _16285_ (.A(_13303_),
    .Y(_13401_));
 sky130_fd_sc_hd__o41ai_1 _16286_ (.A1(_13340_),
    .A2(_13264_),
    .A3(_13265_),
    .A4(_13302_),
    .B1(_13383_),
    .Y(_13402_));
 sky130_fd_sc_hd__a21oi_1 _16287_ (.A1(_13340_),
    .A2(_13401_),
    .B1(_13402_),
    .Y(_03904_));
 sky130_fd_sc_hd__a41oi_1 _16288_ (.A1(\count_instr[37] ),
    .A2(_13301_),
    .A3(\count_instr[36] ),
    .A4(\count_instr[35] ),
    .B1(\count_instr[38] ),
    .Y(_13403_));
 sky130_fd_sc_hd__nor3_1 _16289_ (.A(_13392_),
    .B(_13403_),
    .C(_13303_),
    .Y(_03903_));
 sky130_fd_sc_hd__o21bai_1 _16290_ (.A1(_13265_),
    .A2(_13302_),
    .B1_N(_13386_),
    .Y(_13404_));
 sky130_fd_sc_hd__a21oi_1 _16291_ (.A1(_13265_),
    .A2(_13302_),
    .B1(_13404_),
    .Y(_03902_));
 sky130_fd_sc_hd__a31oi_1 _16292_ (.A1(_13301_),
    .A2(\count_instr[36] ),
    .A3(\count_instr[35] ),
    .B1(_13388_),
    .Y(_13405_));
 sky130_fd_sc_hd__o21a_1 _16293_ (.A1(\count_instr[36] ),
    .A2(_13365_),
    .B1(_13405_),
    .X(_03901_));
 sky130_vsdinv _16294_ (.A(_13301_),
    .Y(_13406_));
 sky130_fd_sc_hd__o41ai_1 _16295_ (.A1(_13341_),
    .A2(_13266_),
    .A3(_13267_),
    .A4(_13300_),
    .B1(_13383_),
    .Y(_13407_));
 sky130_fd_sc_hd__a21oi_1 _16296_ (.A1(_13341_),
    .A2(_13406_),
    .B1(_13407_),
    .Y(_03900_));
 sky130_fd_sc_hd__o31ai_1 _16297_ (.A1(_13266_),
    .A2(_13267_),
    .A3(_13300_),
    .B1(_13333_),
    .Y(_13408_));
 sky130_fd_sc_hd__a21oi_1 _16298_ (.A1(_13266_),
    .A2(_13364_),
    .B1(_13408_),
    .Y(_03899_));
 sky130_fd_sc_hd__o21bai_1 _16299_ (.A1(_13267_),
    .A2(_13300_),
    .B1_N(_13386_),
    .Y(_13409_));
 sky130_fd_sc_hd__a21oi_1 _16300_ (.A1(_13267_),
    .A2(_13300_),
    .B1(_13409_),
    .Y(_03898_));
 sky130_fd_sc_hd__a31oi_1 _16301_ (.A1(_13299_),
    .A2(\count_instr[32] ),
    .A3(\count_instr[31] ),
    .B1(_13388_),
    .Y(_13410_));
 sky130_fd_sc_hd__o21a_1 _16302_ (.A1(\count_instr[32] ),
    .A2(_13363_),
    .B1(_13410_),
    .X(_03897_));
 sky130_vsdinv _16303_ (.A(_13299_),
    .Y(_13411_));
 sky130_fd_sc_hd__o41ai_1 _16304_ (.A1(_13342_),
    .A2(_13268_),
    .A3(_13269_),
    .A4(_13298_),
    .B1(_13383_),
    .Y(_13412_));
 sky130_fd_sc_hd__a21oi_1 _16305_ (.A1(_13342_),
    .A2(_13411_),
    .B1(_13412_),
    .Y(_03896_));
 sky130_fd_sc_hd__a41oi_2 _16306_ (.A1(\count_instr[29] ),
    .A2(_13297_),
    .A3(\count_instr[28] ),
    .A4(\count_instr[27] ),
    .B1(\count_instr[30] ),
    .Y(_13413_));
 sky130_fd_sc_hd__nor3_1 _16307_ (.A(_13392_),
    .B(_13413_),
    .C(_13299_),
    .Y(_03895_));
 sky130_fd_sc_hd__o21bai_1 _16308_ (.A1(_13269_),
    .A2(_13298_),
    .B1_N(_13386_),
    .Y(_13414_));
 sky130_fd_sc_hd__a21oi_1 _16309_ (.A1(_13269_),
    .A2(_13298_),
    .B1(_13414_),
    .Y(_03894_));
 sky130_fd_sc_hd__a31oi_1 _16310_ (.A1(_13297_),
    .A2(\count_instr[28] ),
    .A3(\count_instr[27] ),
    .B1(_13388_),
    .Y(_13415_));
 sky130_fd_sc_hd__o21a_1 _16311_ (.A1(\count_instr[28] ),
    .A2(_13361_),
    .B1(_13415_),
    .X(_03893_));
 sky130_vsdinv _16312_ (.A(_13297_),
    .Y(_13416_));
 sky130_fd_sc_hd__buf_2 _16313_ (.A(_12895_),
    .X(_13417_));
 sky130_fd_sc_hd__o41ai_1 _16314_ (.A1(_13343_),
    .A2(_13270_),
    .A3(_13271_),
    .A4(_13296_),
    .B1(_13417_),
    .Y(_13418_));
 sky130_fd_sc_hd__a21oi_1 _16315_ (.A1(_13343_),
    .A2(_13416_),
    .B1(_13418_),
    .Y(_03892_));
 sky130_fd_sc_hd__o31ai_1 _16316_ (.A1(_13270_),
    .A2(_13271_),
    .A3(_13296_),
    .B1(_13333_),
    .Y(_13419_));
 sky130_fd_sc_hd__a21oi_1 _16317_ (.A1(_13270_),
    .A2(_13360_),
    .B1(_13419_),
    .Y(_03891_));
 sky130_fd_sc_hd__buf_2 _16318_ (.A(_12643_),
    .X(_13420_));
 sky130_fd_sc_hd__o21bai_1 _16319_ (.A1(_13271_),
    .A2(_13296_),
    .B1_N(_13420_),
    .Y(_13421_));
 sky130_fd_sc_hd__a21oi_1 _16320_ (.A1(_13271_),
    .A2(_13296_),
    .B1(_13421_),
    .Y(_03890_));
 sky130_fd_sc_hd__buf_2 _16321_ (.A(_12912_),
    .X(_13422_));
 sky130_fd_sc_hd__a31oi_1 _16322_ (.A1(_13295_),
    .A2(\count_instr[24] ),
    .A3(\count_instr[23] ),
    .B1(_13422_),
    .Y(_13423_));
 sky130_fd_sc_hd__o21a_1 _16323_ (.A1(\count_instr[24] ),
    .A2(_13359_),
    .B1(_13423_),
    .X(_03889_));
 sky130_vsdinv _16324_ (.A(_13295_),
    .Y(_13424_));
 sky130_fd_sc_hd__o41ai_1 _16325_ (.A1(_13344_),
    .A2(_13272_),
    .A3(_13273_),
    .A4(_13294_),
    .B1(_13417_),
    .Y(_13425_));
 sky130_fd_sc_hd__a21oi_1 _16326_ (.A1(_13344_),
    .A2(_13424_),
    .B1(_13425_),
    .Y(_03888_));
 sky130_fd_sc_hd__o31ai_1 _16327_ (.A1(_13272_),
    .A2(_13273_),
    .A3(_13294_),
    .B1(_13333_),
    .Y(_13426_));
 sky130_fd_sc_hd__a21oi_1 _16328_ (.A1(_13272_),
    .A2(_13358_),
    .B1(_13426_),
    .Y(_03887_));
 sky130_fd_sc_hd__o21bai_1 _16329_ (.A1(_13273_),
    .A2(_13294_),
    .B1_N(_13420_),
    .Y(_13427_));
 sky130_fd_sc_hd__a21oi_1 _16330_ (.A1(_13273_),
    .A2(_13294_),
    .B1(_13427_),
    .Y(_03886_));
 sky130_fd_sc_hd__a31oi_1 _16331_ (.A1(_13293_),
    .A2(\count_instr[20] ),
    .A3(\count_instr[19] ),
    .B1(_13422_),
    .Y(_13428_));
 sky130_fd_sc_hd__o21a_1 _16332_ (.A1(\count_instr[20] ),
    .A2(_13357_),
    .B1(_13428_),
    .X(_03885_));
 sky130_vsdinv _16333_ (.A(_13293_),
    .Y(_13429_));
 sky130_fd_sc_hd__o41ai_1 _16334_ (.A1(_13345_),
    .A2(_13274_),
    .A3(_13275_),
    .A4(_13292_),
    .B1(_13417_),
    .Y(_13430_));
 sky130_fd_sc_hd__a21oi_1 _16335_ (.A1(_13345_),
    .A2(_13429_),
    .B1(_13430_),
    .Y(_03884_));
 sky130_fd_sc_hd__o31ai_1 _16336_ (.A1(_13274_),
    .A2(_13275_),
    .A3(_13292_),
    .B1(_13333_),
    .Y(_13431_));
 sky130_fd_sc_hd__a21oi_1 _16337_ (.A1(_13274_),
    .A2(_13356_),
    .B1(_13431_),
    .Y(_03883_));
 sky130_fd_sc_hd__o21bai_1 _16338_ (.A1(_13275_),
    .A2(_13292_),
    .B1_N(_13420_),
    .Y(_13432_));
 sky130_fd_sc_hd__a21oi_1 _16339_ (.A1(_13275_),
    .A2(_13292_),
    .B1(_13432_),
    .Y(_03882_));
 sky130_fd_sc_hd__a31oi_1 _16340_ (.A1(_13291_),
    .A2(\count_instr[16] ),
    .A3(\count_instr[15] ),
    .B1(_13422_),
    .Y(_13433_));
 sky130_fd_sc_hd__o21a_1 _16341_ (.A1(\count_instr[16] ),
    .A2(_13355_),
    .B1(_13433_),
    .X(_03881_));
 sky130_vsdinv _16342_ (.A(_13291_),
    .Y(_13434_));
 sky130_fd_sc_hd__o41ai_1 _16343_ (.A1(_13346_),
    .A2(_13276_),
    .A3(_13277_),
    .A4(_13290_),
    .B1(_13417_),
    .Y(_13435_));
 sky130_fd_sc_hd__a21oi_1 _16344_ (.A1(_13346_),
    .A2(_13434_),
    .B1(_13435_),
    .Y(_03880_));
 sky130_fd_sc_hd__a41oi_1 _16345_ (.A1(\count_instr[13] ),
    .A2(_13289_),
    .A3(\count_instr[12] ),
    .A4(\count_instr[11] ),
    .B1(\count_instr[14] ),
    .Y(_13436_));
 sky130_fd_sc_hd__nor3_1 _16346_ (.A(_13392_),
    .B(_13436_),
    .C(_13291_),
    .Y(_03879_));
 sky130_fd_sc_hd__o21bai_1 _16347_ (.A1(_13277_),
    .A2(_13290_),
    .B1_N(_13420_),
    .Y(_13437_));
 sky130_fd_sc_hd__a21oi_1 _16348_ (.A1(_13277_),
    .A2(_13290_),
    .B1(_13437_),
    .Y(_03878_));
 sky130_fd_sc_hd__a31oi_1 _16349_ (.A1(_13289_),
    .A2(\count_instr[12] ),
    .A3(\count_instr[11] ),
    .B1(_13422_),
    .Y(_13438_));
 sky130_fd_sc_hd__o21a_1 _16350_ (.A1(\count_instr[12] ),
    .A2(_13353_),
    .B1(_13438_),
    .X(_03877_));
 sky130_vsdinv _16351_ (.A(_13289_),
    .Y(_13439_));
 sky130_fd_sc_hd__o41ai_1 _16352_ (.A1(_13347_),
    .A2(_13278_),
    .A3(_13279_),
    .A4(_13288_),
    .B1(_13417_),
    .Y(_13440_));
 sky130_fd_sc_hd__a21oi_1 _16353_ (.A1(_13347_),
    .A2(_13439_),
    .B1(_13440_),
    .Y(_03876_));
 sky130_fd_sc_hd__a41oi_1 _16354_ (.A1(\count_instr[9] ),
    .A2(_13287_),
    .A3(\count_instr[8] ),
    .A4(\count_instr[7] ),
    .B1(\count_instr[10] ),
    .Y(_13441_));
 sky130_fd_sc_hd__nor3_1 _16355_ (.A(_13392_),
    .B(_13441_),
    .C(_13289_),
    .Y(_03875_));
 sky130_fd_sc_hd__o21bai_1 _16356_ (.A1(_13279_),
    .A2(_13288_),
    .B1_N(_13420_),
    .Y(_13442_));
 sky130_fd_sc_hd__a21oi_1 _16357_ (.A1(_13279_),
    .A2(_13288_),
    .B1(_13442_),
    .Y(_03874_));
 sky130_fd_sc_hd__a31oi_1 _16358_ (.A1(_13287_),
    .A2(\count_instr[8] ),
    .A3(\count_instr[7] ),
    .B1(_13422_),
    .Y(_13443_));
 sky130_fd_sc_hd__o21a_1 _16359_ (.A1(\count_instr[8] ),
    .A2(_13351_),
    .B1(_13443_),
    .X(_03873_));
 sky130_vsdinv _16360_ (.A(_13287_),
    .Y(_13444_));
 sky130_fd_sc_hd__o41ai_1 _16361_ (.A1(_13348_),
    .A2(_13280_),
    .A3(_13281_),
    .A4(_13286_),
    .B1(_13417_),
    .Y(_13445_));
 sky130_fd_sc_hd__a21oi_1 _16362_ (.A1(_13348_),
    .A2(_13444_),
    .B1(_13445_),
    .Y(_03872_));
 sky130_fd_sc_hd__o31ai_1 _16363_ (.A1(_13280_),
    .A2(_13281_),
    .A3(_13286_),
    .B1(_12920_),
    .Y(_13446_));
 sky130_fd_sc_hd__a21oi_1 _16364_ (.A1(_13280_),
    .A2(_13350_),
    .B1(_13446_),
    .Y(_03871_));
 sky130_fd_sc_hd__o21bai_1 _16365_ (.A1(_13281_),
    .A2(_13286_),
    .B1_N(_13420_),
    .Y(_13447_));
 sky130_fd_sc_hd__a21oi_1 _16366_ (.A1(_13281_),
    .A2(_13286_),
    .B1(_13447_),
    .Y(_03870_));
 sky130_fd_sc_hd__a31oi_1 _16367_ (.A1(_13285_),
    .A2(\count_instr[4] ),
    .A3(\count_instr[3] ),
    .B1(_13422_),
    .Y(_13448_));
 sky130_fd_sc_hd__o21a_1 _16368_ (.A1(\count_instr[4] ),
    .A2(_13349_),
    .B1(_13448_),
    .X(_03869_));
 sky130_fd_sc_hd__a21oi_1 _16369_ (.A1(_13285_),
    .A2(\count_instr[3] ),
    .B1(_12964_),
    .Y(_13449_));
 sky130_fd_sc_hd__o21a_1 _16370_ (.A1(\count_instr[3] ),
    .A2(_13285_),
    .B1(_13449_),
    .X(_03868_));
 sky130_fd_sc_hd__nor3b_4 _16371_ (.A(_13282_),
    .B(_12901_),
    .C_N(\count_instr[1] ),
    .Y(_13450_));
 sky130_vsdinv _16372_ (.A(_13285_),
    .Y(_13451_));
 sky130_fd_sc_hd__o211a_1 _16373_ (.A1(\count_instr[2] ),
    .A2(_13450_),
    .B1(_13238_),
    .C1(_13451_),
    .X(_03867_));
 sky130_fd_sc_hd__clkbuf_4 _16374_ (.A(_13321_),
    .X(_13452_));
 sky130_fd_sc_hd__o21ba_1 _16375_ (.A1(_13282_),
    .A2(_12901_),
    .B1_N(\count_instr[1] ),
    .X(_13453_));
 sky130_fd_sc_hd__nor3_1 _16376_ (.A(_13452_),
    .B(_13450_),
    .C(_13453_),
    .Y(_03866_));
 sky130_fd_sc_hd__o21bai_1 _16377_ (.A1(_13282_),
    .A2(_12901_),
    .B1_N(_12912_),
    .Y(_13454_));
 sky130_fd_sc_hd__a21oi_1 _16378_ (.A1(_13282_),
    .A2(_12901_),
    .B1(_13454_),
    .Y(_03865_));
 sky130_fd_sc_hd__inv_2 _16379_ (.A(_12861_),
    .Y(_13455_));
 sky130_fd_sc_hd__nor2_2 _16380_ (.A(\cpu_state[1] ),
    .B(\cpu_state[2] ),
    .Y(_00315_));
 sky130_fd_sc_hd__a211o_2 _16381_ (.A1(_13455_),
    .A2(\cpu_state[1] ),
    .B1(_00315_),
    .C1(_12662_),
    .X(_13456_));
 sky130_fd_sc_hd__buf_2 _16382_ (.A(_13456_),
    .X(_13457_));
 sky130_fd_sc_hd__clkbuf_2 _16383_ (.A(_13457_),
    .X(_13458_));
 sky130_fd_sc_hd__clkbuf_4 _16384_ (.A(_12916_),
    .X(_13459_));
 sky130_fd_sc_hd__nor3b_1 _16385_ (.A(\irq_mask[31] ),
    .B(_13459_),
    .C_N(\irq_pending[31] ),
    .Y(_13460_));
 sky130_fd_sc_hd__clkbuf_2 _16386_ (.A(_13195_),
    .X(_13461_));
 sky130_fd_sc_hd__clkbuf_2 _16387_ (.A(_13456_),
    .X(_13462_));
 sky130_fd_sc_hd__or2b_1 _16388_ (.A(net126),
    .B_N(_13462_),
    .X(_13463_));
 sky130_fd_sc_hd__o211a_1 _16389_ (.A1(_13458_),
    .A2(_13460_),
    .B1(_13461_),
    .C1(_13463_),
    .X(_03864_));
 sky130_fd_sc_hd__nor3b_2 _16390_ (.A(\irq_mask[30] ),
    .B(_13459_),
    .C_N(\irq_pending[30] ),
    .Y(_13464_));
 sky130_fd_sc_hd__or2b_1 _16391_ (.A(net125),
    .B_N(_13462_),
    .X(_13465_));
 sky130_fd_sc_hd__o211a_1 _16392_ (.A1(_13458_),
    .A2(_13464_),
    .B1(_13461_),
    .C1(_13465_),
    .X(_03863_));
 sky130_fd_sc_hd__nor3b_2 _16393_ (.A(\irq_mask[29] ),
    .B(_13459_),
    .C_N(\irq_pending[29] ),
    .Y(_13466_));
 sky130_fd_sc_hd__or2b_1 _16394_ (.A(net123),
    .B_N(_13462_),
    .X(_13467_));
 sky130_fd_sc_hd__o211a_1 _16395_ (.A1(_13458_),
    .A2(_13466_),
    .B1(_13461_),
    .C1(_13467_),
    .X(_03862_));
 sky130_fd_sc_hd__nor3b_2 _16396_ (.A(\irq_mask[28] ),
    .B(_13459_),
    .C_N(\irq_pending[28] ),
    .Y(_13468_));
 sky130_fd_sc_hd__or2b_1 _16397_ (.A(net122),
    .B_N(_13462_),
    .X(_13469_));
 sky130_fd_sc_hd__o211a_1 _16398_ (.A1(_13458_),
    .A2(_13468_),
    .B1(_13461_),
    .C1(_13469_),
    .X(_03861_));
 sky130_fd_sc_hd__nor3b_2 _16399_ (.A(\irq_mask[27] ),
    .B(_13459_),
    .C_N(\irq_pending[27] ),
    .Y(_13470_));
 sky130_fd_sc_hd__clkbuf_2 _16400_ (.A(_13456_),
    .X(_13471_));
 sky130_fd_sc_hd__buf_2 _16401_ (.A(_13471_),
    .X(_13472_));
 sky130_fd_sc_hd__or2b_1 _16402_ (.A(net121),
    .B_N(_13472_),
    .X(_13473_));
 sky130_fd_sc_hd__o211a_1 _16403_ (.A1(_13458_),
    .A2(_13470_),
    .B1(_13461_),
    .C1(_13473_),
    .X(_03860_));
 sky130_fd_sc_hd__nor3b_2 _16404_ (.A(\irq_mask[26] ),
    .B(_13459_),
    .C_N(\irq_pending[26] ),
    .Y(_13474_));
 sky130_fd_sc_hd__or2b_1 _16405_ (.A(net120),
    .B_N(_13472_),
    .X(_13475_));
 sky130_fd_sc_hd__o211a_1 _16406_ (.A1(_13458_),
    .A2(_13474_),
    .B1(_13461_),
    .C1(_13475_),
    .X(_03859_));
 sky130_fd_sc_hd__buf_2 _16407_ (.A(_13457_),
    .X(_13476_));
 sky130_fd_sc_hd__clkbuf_4 _16408_ (.A(_12915_),
    .X(_13477_));
 sky130_fd_sc_hd__nor3b_2 _16409_ (.A(\irq_mask[25] ),
    .B(_13477_),
    .C_N(\irq_pending[25] ),
    .Y(_13478_));
 sky130_fd_sc_hd__buf_2 _16410_ (.A(_13195_),
    .X(_13479_));
 sky130_fd_sc_hd__or2b_1 _16411_ (.A(net119),
    .B_N(_13472_),
    .X(_13480_));
 sky130_fd_sc_hd__o211a_1 _16412_ (.A1(_13476_),
    .A2(_13478_),
    .B1(_13479_),
    .C1(_13480_),
    .X(_03858_));
 sky130_fd_sc_hd__nor3b_2 _16413_ (.A(\irq_mask[24] ),
    .B(_13477_),
    .C_N(\irq_pending[24] ),
    .Y(_13481_));
 sky130_fd_sc_hd__or2b_1 _16414_ (.A(net118),
    .B_N(_13472_),
    .X(_13482_));
 sky130_fd_sc_hd__o211a_1 _16415_ (.A1(_13476_),
    .A2(_13481_),
    .B1(_13479_),
    .C1(_13482_),
    .X(_03857_));
 sky130_fd_sc_hd__nor3b_1 _16416_ (.A(\irq_mask[23] ),
    .B(_13477_),
    .C_N(\irq_pending[23] ),
    .Y(_13483_));
 sky130_fd_sc_hd__or2b_1 _16417_ (.A(net117),
    .B_N(_13472_),
    .X(_13484_));
 sky130_fd_sc_hd__o211a_1 _16418_ (.A1(_13476_),
    .A2(_13483_),
    .B1(_13479_),
    .C1(_13484_),
    .X(_03856_));
 sky130_fd_sc_hd__nor3b_2 _16419_ (.A(\irq_mask[22] ),
    .B(_13477_),
    .C_N(\irq_pending[22] ),
    .Y(_13485_));
 sky130_fd_sc_hd__or2b_1 _16420_ (.A(net116),
    .B_N(_13472_),
    .X(_13486_));
 sky130_fd_sc_hd__o211a_1 _16421_ (.A1(_13476_),
    .A2(_13485_),
    .B1(_13479_),
    .C1(_13486_),
    .X(_03855_));
 sky130_fd_sc_hd__nor3b_1 _16422_ (.A(\irq_mask[21] ),
    .B(_13477_),
    .C_N(\irq_pending[21] ),
    .Y(_13487_));
 sky130_fd_sc_hd__clkbuf_2 _16423_ (.A(_13471_),
    .X(_13488_));
 sky130_fd_sc_hd__or2b_1 _16424_ (.A(net115),
    .B_N(_13488_),
    .X(_13489_));
 sky130_fd_sc_hd__o211a_1 _16425_ (.A1(_13476_),
    .A2(_13487_),
    .B1(_13479_),
    .C1(_13489_),
    .X(_03854_));
 sky130_fd_sc_hd__nor3b_2 _16426_ (.A(\irq_mask[20] ),
    .B(_13477_),
    .C_N(\irq_pending[20] ),
    .Y(_13490_));
 sky130_fd_sc_hd__or2b_1 _16427_ (.A(net114),
    .B_N(_13488_),
    .X(_13491_));
 sky130_fd_sc_hd__o211a_1 _16428_ (.A1(_13476_),
    .A2(_13490_),
    .B1(_13479_),
    .C1(_13491_),
    .X(_03853_));
 sky130_fd_sc_hd__clkbuf_2 _16429_ (.A(_13471_),
    .X(_13492_));
 sky130_fd_sc_hd__clkbuf_4 _16430_ (.A(_12915_),
    .X(_13493_));
 sky130_fd_sc_hd__nor3b_2 _16431_ (.A(\irq_mask[19] ),
    .B(_13493_),
    .C_N(\irq_pending[19] ),
    .Y(_13494_));
 sky130_fd_sc_hd__clkbuf_2 _16432_ (.A(_13195_),
    .X(_13495_));
 sky130_fd_sc_hd__or2b_1 _16433_ (.A(net112),
    .B_N(_13488_),
    .X(_13496_));
 sky130_fd_sc_hd__o211a_1 _16434_ (.A1(_13492_),
    .A2(_13494_),
    .B1(_13495_),
    .C1(_13496_),
    .X(_03852_));
 sky130_fd_sc_hd__nor3b_1 _16435_ (.A(\irq_mask[18] ),
    .B(_13493_),
    .C_N(\irq_pending[18] ),
    .Y(_13497_));
 sky130_fd_sc_hd__or2b_1 _16436_ (.A(net111),
    .B_N(_13488_),
    .X(_13498_));
 sky130_fd_sc_hd__o211a_1 _16437_ (.A1(_13492_),
    .A2(_13497_),
    .B1(_13495_),
    .C1(_13498_),
    .X(_03851_));
 sky130_fd_sc_hd__nor3b_1 _16438_ (.A(\irq_mask[17] ),
    .B(_13493_),
    .C_N(\irq_pending[17] ),
    .Y(_13499_));
 sky130_fd_sc_hd__or2b_1 _16439_ (.A(net110),
    .B_N(_13488_),
    .X(_13500_));
 sky130_fd_sc_hd__o211a_1 _16440_ (.A1(_13492_),
    .A2(_13499_),
    .B1(_13495_),
    .C1(_13500_),
    .X(_03850_));
 sky130_fd_sc_hd__nor3b_2 _16441_ (.A(\irq_mask[16] ),
    .B(_13493_),
    .C_N(\irq_pending[16] ),
    .Y(_13501_));
 sky130_fd_sc_hd__or2b_1 _16442_ (.A(net109),
    .B_N(_13488_),
    .X(_13502_));
 sky130_fd_sc_hd__o211a_1 _16443_ (.A1(_13492_),
    .A2(_13501_),
    .B1(_13495_),
    .C1(_13502_),
    .X(_03849_));
 sky130_fd_sc_hd__nor3b_2 _16444_ (.A(\irq_mask[15] ),
    .B(_13493_),
    .C_N(\irq_pending[15] ),
    .Y(_13503_));
 sky130_fd_sc_hd__clkbuf_2 _16445_ (.A(_13471_),
    .X(_13504_));
 sky130_fd_sc_hd__or2b_1 _16446_ (.A(net108),
    .B_N(_13504_),
    .X(_13505_));
 sky130_fd_sc_hd__o211a_1 _16447_ (.A1(_13492_),
    .A2(_13503_),
    .B1(_13495_),
    .C1(_13505_),
    .X(_03848_));
 sky130_fd_sc_hd__nor3b_2 _16448_ (.A(\irq_mask[14] ),
    .B(_13493_),
    .C_N(\irq_pending[14] ),
    .Y(_13506_));
 sky130_fd_sc_hd__or2b_1 _16449_ (.A(net107),
    .B_N(_13504_),
    .X(_13507_));
 sky130_fd_sc_hd__o211a_1 _16450_ (.A1(_13492_),
    .A2(_13506_),
    .B1(_13495_),
    .C1(_13507_),
    .X(_03847_));
 sky130_fd_sc_hd__clkbuf_2 _16451_ (.A(_13471_),
    .X(_13508_));
 sky130_fd_sc_hd__clkbuf_4 _16452_ (.A(_12915_),
    .X(_13509_));
 sky130_fd_sc_hd__nor3b_2 _16453_ (.A(\irq_mask[13] ),
    .B(_13509_),
    .C_N(\irq_pending[13] ),
    .Y(_13510_));
 sky130_fd_sc_hd__clkbuf_2 _16454_ (.A(_12649_),
    .X(_13511_));
 sky130_fd_sc_hd__or2b_1 _16455_ (.A(net106),
    .B_N(_13504_),
    .X(_13512_));
 sky130_fd_sc_hd__o211a_1 _16456_ (.A1(_13508_),
    .A2(_13510_),
    .B1(_13511_),
    .C1(_13512_),
    .X(_03846_));
 sky130_fd_sc_hd__nor3b_2 _16457_ (.A(\irq_mask[12] ),
    .B(_13509_),
    .C_N(\irq_pending[12] ),
    .Y(_13513_));
 sky130_fd_sc_hd__or2b_1 _16458_ (.A(net105),
    .B_N(_13504_),
    .X(_13514_));
 sky130_fd_sc_hd__o211a_1 _16459_ (.A1(_13508_),
    .A2(_13513_),
    .B1(_13511_),
    .C1(_13514_),
    .X(_03845_));
 sky130_fd_sc_hd__nor3b_2 _16460_ (.A(\irq_mask[11] ),
    .B(_13509_),
    .C_N(\irq_pending[11] ),
    .Y(_13515_));
 sky130_fd_sc_hd__or2b_1 _16461_ (.A(net104),
    .B_N(_13504_),
    .X(_13516_));
 sky130_fd_sc_hd__o211a_1 _16462_ (.A1(_13508_),
    .A2(_13515_),
    .B1(_13511_),
    .C1(_13516_),
    .X(_03844_));
 sky130_fd_sc_hd__nor3b_2 _16463_ (.A(\irq_mask[10] ),
    .B(_13509_),
    .C_N(\irq_pending[10] ),
    .Y(_13517_));
 sky130_fd_sc_hd__or2b_1 _16464_ (.A(net103),
    .B_N(_13504_),
    .X(_13518_));
 sky130_fd_sc_hd__o211a_1 _16465_ (.A1(_13508_),
    .A2(_13517_),
    .B1(_13511_),
    .C1(_13518_),
    .X(_03843_));
 sky130_fd_sc_hd__nor3b_2 _16466_ (.A(\irq_mask[9] ),
    .B(_13509_),
    .C_N(\irq_pending[9] ),
    .Y(_13519_));
 sky130_fd_sc_hd__clkbuf_2 _16467_ (.A(_13456_),
    .X(_13520_));
 sky130_fd_sc_hd__or2b_1 _16468_ (.A(net133),
    .B_N(_13520_),
    .X(_13521_));
 sky130_fd_sc_hd__o211a_1 _16469_ (.A1(_13508_),
    .A2(_13519_),
    .B1(_13511_),
    .C1(_13521_),
    .X(_03842_));
 sky130_fd_sc_hd__nor3b_2 _16470_ (.A(\irq_mask[8] ),
    .B(_13509_),
    .C_N(\irq_pending[8] ),
    .Y(_13522_));
 sky130_fd_sc_hd__or2b_1 _16471_ (.A(net132),
    .B_N(_13520_),
    .X(_13523_));
 sky130_fd_sc_hd__o211a_1 _16472_ (.A1(_13508_),
    .A2(_13522_),
    .B1(_13511_),
    .C1(_13523_),
    .X(_03841_));
 sky130_fd_sc_hd__clkbuf_2 _16473_ (.A(_13471_),
    .X(_13524_));
 sky130_fd_sc_hd__buf_2 _16474_ (.A(_12915_),
    .X(_13525_));
 sky130_fd_sc_hd__nor3b_1 _16475_ (.A(\irq_mask[7] ),
    .B(_13525_),
    .C_N(\irq_pending[7] ),
    .Y(_13526_));
 sky130_fd_sc_hd__clkbuf_2 _16476_ (.A(_12649_),
    .X(_13527_));
 sky130_fd_sc_hd__or2b_1 _16477_ (.A(net131),
    .B_N(_13520_),
    .X(_13528_));
 sky130_fd_sc_hd__o211a_1 _16478_ (.A1(_13524_),
    .A2(_13526_),
    .B1(_13527_),
    .C1(_13528_),
    .X(_03840_));
 sky130_fd_sc_hd__nor3b_2 _16479_ (.A(\irq_mask[6] ),
    .B(_13525_),
    .C_N(\irq_pending[6] ),
    .Y(_13529_));
 sky130_fd_sc_hd__or2b_1 _16480_ (.A(net130),
    .B_N(_13520_),
    .X(_13530_));
 sky130_fd_sc_hd__o211a_1 _16481_ (.A1(_13524_),
    .A2(_13529_),
    .B1(_13527_),
    .C1(_13530_),
    .X(_03839_));
 sky130_fd_sc_hd__nor3b_2 _16482_ (.A(\irq_mask[5] ),
    .B(_13525_),
    .C_N(\irq_pending[5] ),
    .Y(_13531_));
 sky130_fd_sc_hd__or2b_1 _16483_ (.A(net129),
    .B_N(_13520_),
    .X(_13532_));
 sky130_fd_sc_hd__o211a_1 _16484_ (.A1(_13524_),
    .A2(_13531_),
    .B1(_13527_),
    .C1(_13532_),
    .X(_03838_));
 sky130_fd_sc_hd__nor3b_2 _16485_ (.A(\irq_mask[4] ),
    .B(_13525_),
    .C_N(\irq_pending[4] ),
    .Y(_13533_));
 sky130_fd_sc_hd__or2b_1 _16486_ (.A(net128),
    .B_N(_13520_),
    .X(_13534_));
 sky130_fd_sc_hd__o211a_1 _16487_ (.A1(_13524_),
    .A2(_13533_),
    .B1(_13527_),
    .C1(_13534_),
    .X(_03837_));
 sky130_fd_sc_hd__nor3b_2 _16488_ (.A(\irq_mask[3] ),
    .B(_13525_),
    .C_N(\irq_pending[3] ),
    .Y(_13535_));
 sky130_fd_sc_hd__or2b_1 _16489_ (.A(net127),
    .B_N(_13457_),
    .X(_13536_));
 sky130_fd_sc_hd__o211a_1 _16490_ (.A1(_13524_),
    .A2(_13535_),
    .B1(_13527_),
    .C1(_13536_),
    .X(_03836_));
 sky130_fd_sc_hd__buf_2 _16491_ (.A(\irq_mask[2] ),
    .X(_13537_));
 sky130_fd_sc_hd__nor3b_2 _16492_ (.A(_13537_),
    .B(_13525_),
    .C_N(\irq_pending[2] ),
    .Y(_13538_));
 sky130_fd_sc_hd__or2b_1 _16493_ (.A(net124),
    .B_N(_13457_),
    .X(_13539_));
 sky130_fd_sc_hd__o211a_1 _16494_ (.A1(_13524_),
    .A2(_13538_),
    .B1(_13527_),
    .C1(_13539_),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_4 _16495_ (.A(\irq_mask[1] ),
    .X(_13540_));
 sky130_fd_sc_hd__nor3b_4 _16496_ (.A(_13540_),
    .B(_12916_),
    .C_N(\irq_pending[1] ),
    .Y(_13541_));
 sky130_fd_sc_hd__buf_4 _16497_ (.A(_12649_),
    .X(_13542_));
 sky130_fd_sc_hd__or2b_1 _16498_ (.A(net113),
    .B_N(_13457_),
    .X(_13543_));
 sky130_fd_sc_hd__o211a_1 _16499_ (.A1(_13462_),
    .A2(_13541_),
    .B1(_13542_),
    .C1(_13543_),
    .X(_03834_));
 sky130_fd_sc_hd__nor3b_4 _16500_ (.A(\irq_mask[0] ),
    .B(_12916_),
    .C_N(\irq_pending[0] ),
    .Y(_13544_));
 sky130_fd_sc_hd__or2b_1 _16501_ (.A(net102),
    .B_N(_13457_),
    .X(_13545_));
 sky130_fd_sc_hd__o211a_1 _16502_ (.A1(_13462_),
    .A2(_13544_),
    .B1(_13542_),
    .C1(_13545_),
    .X(_03833_));
 sky130_fd_sc_hd__and3_1 _16503_ (.A(_12886_),
    .B(_12842_),
    .C(_12887_),
    .X(_13546_));
 sky130_fd_sc_hd__nor2_2 _16504_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_00311_));
 sky130_vsdinv _16505_ (.A(_00311_),
    .Y(_13547_));
 sky130_fd_sc_hd__buf_6 _16506_ (.A(_12885_),
    .X(_13548_));
 sky130_fd_sc_hd__o2111ai_2 _16507_ (.A1(\pcpi_mul.active[1] ),
    .A2(_13547_),
    .B1(_13548_),
    .C1(_12887_),
    .D1(_12886_),
    .Y(_13549_));
 sky130_fd_sc_hd__o211a_1 _16508_ (.A1(net370),
    .A2(_13546_),
    .B1(_13542_),
    .C1(_13549_),
    .X(_03832_));
 sky130_fd_sc_hd__o21a_1 _16509_ (.A1(_00290_),
    .A2(_12630_),
    .B1(net237),
    .X(_13550_));
 sky130_fd_sc_hd__o21bai_1 _16510_ (.A1(_12973_),
    .A2(_13550_),
    .B1_N(net408),
    .Y(_13551_));
 sky130_fd_sc_hd__nand2_1 _16511_ (.A(_12634_),
    .B(net237),
    .Y(_13552_));
 sky130_fd_sc_hd__a21oi_1 _16512_ (.A1(_13551_),
    .A2(_13552_),
    .B1(_13322_),
    .Y(_03831_));
 sky130_fd_sc_hd__or4_4 _16513_ (.A(\irq_pending[25] ),
    .B(\irq_pending[24] ),
    .C(\irq_pending[27] ),
    .D(\irq_pending[26] ),
    .X(_13553_));
 sky130_fd_sc_hd__or4_4 _16514_ (.A(\irq_pending[21] ),
    .B(\irq_pending[20] ),
    .C(\irq_pending[23] ),
    .D(\irq_pending[22] ),
    .X(_13554_));
 sky130_fd_sc_hd__or4_4 _16515_ (.A(\irq_pending[17] ),
    .B(\irq_pending[16] ),
    .C(\irq_pending[19] ),
    .D(\irq_pending[18] ),
    .X(_13555_));
 sky130_fd_sc_hd__or4_4 _16516_ (.A(\irq_pending[29] ),
    .B(\irq_pending[28] ),
    .C(\irq_pending[31] ),
    .D(\irq_pending[30] ),
    .X(_13556_));
 sky130_fd_sc_hd__nor3_2 _16517_ (.A(_13554_),
    .B(_13555_),
    .C(_13556_),
    .Y(_13557_));
 sky130_fd_sc_hd__or2b_4 _16518_ (.A(_13553_),
    .B_N(_13557_),
    .X(_13558_));
 sky130_fd_sc_hd__or4_4 _16519_ (.A(\irq_pending[9] ),
    .B(\irq_pending[8] ),
    .C(\irq_pending[11] ),
    .D(\irq_pending[10] ),
    .X(_13559_));
 sky130_fd_sc_hd__or4_4 _16520_ (.A(\irq_pending[5] ),
    .B(\irq_pending[4] ),
    .C(\irq_pending[7] ),
    .D(\irq_pending[6] ),
    .X(_13560_));
 sky130_fd_sc_hd__or4_4 _16521_ (.A(\irq_pending[1] ),
    .B(\irq_pending[0] ),
    .C(\irq_pending[3] ),
    .D(\irq_pending[2] ),
    .X(_13561_));
 sky130_fd_sc_hd__or4_4 _16522_ (.A(\irq_pending[13] ),
    .B(\irq_pending[12] ),
    .C(\irq_pending[15] ),
    .D(\irq_pending[14] ),
    .X(_13562_));
 sky130_fd_sc_hd__nor3_2 _16523_ (.A(_13560_),
    .B(_13561_),
    .C(_13562_),
    .Y(_13563_));
 sky130_fd_sc_hd__or2b_2 _16524_ (.A(_13559_),
    .B_N(_13563_),
    .X(_13564_));
 sky130_fd_sc_hd__nor2_4 _16525_ (.A(_13558_),
    .B(_13564_),
    .Y(_02410_));
 sky130_vsdinv _16526_ (.A(_00309_),
    .Y(_13565_));
 sky130_fd_sc_hd__nand3_4 _16527_ (.A(_12771_),
    .B(net101),
    .C(_12873_),
    .Y(_13566_));
 sky130_fd_sc_hd__and2b_1 _16528_ (.A_N(_13559_),
    .B(_13563_),
    .X(_13567_));
 sky130_fd_sc_hd__nand3b_2 _16529_ (.A_N(_13558_),
    .B(_12879_),
    .C(_13567_),
    .Y(_13568_));
 sky130_fd_sc_hd__nor3_1 _16530_ (.A(_13565_),
    .B(_13566_),
    .C(_13568_),
    .Y(_03830_));
 sky130_fd_sc_hd__nor2_4 _16531_ (.A(instr_sltu),
    .B(instr_sltiu),
    .Y(_13569_));
 sky130_fd_sc_hd__nor2_4 _16532_ (.A(instr_slt),
    .B(instr_slti),
    .Y(_13570_));
 sky130_vsdinv _16533_ (.A(_12978_),
    .Y(_13571_));
 sky130_fd_sc_hd__clkbuf_4 _16534_ (.A(_13070_),
    .X(_13572_));
 sky130_fd_sc_hd__a311oi_4 _16535_ (.A1(_13569_),
    .A2(_13570_),
    .A3(_13571_),
    .B1(_13169_),
    .C1(_13572_),
    .Y(_03829_));
 sky130_fd_sc_hd__nand3_4 _16536_ (.A(_12632_),
    .B(net456),
    .C(_13089_),
    .Y(_13573_));
 sky130_fd_sc_hd__nor3_4 _16537_ (.A(_12642_),
    .B(_00297_),
    .C(_13573_),
    .Y(_03828_));
 sky130_fd_sc_hd__nor2_1 _16538_ (.A(_12872_),
    .B(_13087_),
    .Y(_03827_));
 sky130_fd_sc_hd__and2_1 _16539_ (.A(_12971_),
    .B(_02435_),
    .X(_03826_));
 sky130_fd_sc_hd__and2_1 _16540_ (.A(_12971_),
    .B(_02434_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_1 _16541_ (.A(_12971_),
    .B(_02432_),
    .X(_03824_));
 sky130_fd_sc_hd__and2_1 _16542_ (.A(_12971_),
    .B(_02431_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_2 _16543_ (.A(_12961_),
    .X(_13574_));
 sky130_fd_sc_hd__and2_1 _16544_ (.A(_13574_),
    .B(_02430_),
    .X(_03822_));
 sky130_fd_sc_hd__and2_1 _16545_ (.A(_13574_),
    .B(_02429_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_1 _16546_ (.A(_13574_),
    .B(_02428_),
    .X(_03820_));
 sky130_fd_sc_hd__and2_1 _16547_ (.A(_13574_),
    .B(_02427_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_1 _16548_ (.A(_13574_),
    .B(_02426_),
    .X(_03818_));
 sky130_fd_sc_hd__and2_1 _16549_ (.A(_13574_),
    .B(_02425_),
    .X(_03817_));
 sky130_fd_sc_hd__buf_1 _16550_ (.A(_12961_),
    .X(_13575_));
 sky130_fd_sc_hd__and2_1 _16551_ (.A(_13575_),
    .B(_02424_),
    .X(_03816_));
 sky130_fd_sc_hd__and2_1 _16552_ (.A(_13575_),
    .B(_02423_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_1 _16553_ (.A(_13575_),
    .B(_02421_),
    .X(_03814_));
 sky130_fd_sc_hd__and2_1 _16554_ (.A(_13575_),
    .B(_02420_),
    .X(_03813_));
 sky130_fd_sc_hd__and2_1 _16555_ (.A(_13575_),
    .B(_02419_),
    .X(_03812_));
 sky130_fd_sc_hd__and2_1 _16556_ (.A(_13575_),
    .B(_02418_),
    .X(_03811_));
 sky130_fd_sc_hd__clkbuf_2 _16557_ (.A(_12961_),
    .X(_13576_));
 sky130_fd_sc_hd__and2_1 _16558_ (.A(_13576_),
    .B(_02417_),
    .X(_03810_));
 sky130_fd_sc_hd__and2_1 _16559_ (.A(_13576_),
    .B(_02416_),
    .X(_03809_));
 sky130_fd_sc_hd__and2_1 _16560_ (.A(_13576_),
    .B(_02415_),
    .X(_03808_));
 sky130_fd_sc_hd__and2_1 _16561_ (.A(_13576_),
    .B(_02414_),
    .X(_03807_));
 sky130_fd_sc_hd__and2_1 _16562_ (.A(_13576_),
    .B(_02413_),
    .X(_03806_));
 sky130_fd_sc_hd__and2_1 _16563_ (.A(_13576_),
    .B(_02412_),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_2 _16564_ (.A(_12961_),
    .X(_13577_));
 sky130_fd_sc_hd__and2_1 _16565_ (.A(_13577_),
    .B(_02442_),
    .X(_03804_));
 sky130_fd_sc_hd__and2_1 _16566_ (.A(_13577_),
    .B(_02441_),
    .X(_03803_));
 sky130_fd_sc_hd__and2_1 _16567_ (.A(_13577_),
    .B(_02440_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_1 _16568_ (.A(_13577_),
    .B(_02439_),
    .X(_03801_));
 sky130_fd_sc_hd__and2_1 _16569_ (.A(_13577_),
    .B(_02438_),
    .X(_03800_));
 sky130_fd_sc_hd__and2_1 _16570_ (.A(_13577_),
    .B(_02437_),
    .X(_03799_));
 sky130_fd_sc_hd__buf_2 _16571_ (.A(_12961_),
    .X(_13578_));
 sky130_fd_sc_hd__and2_1 _16572_ (.A(_13578_),
    .B(_02436_),
    .X(_03798_));
 sky130_fd_sc_hd__and2_1 _16573_ (.A(_13578_),
    .B(_02433_),
    .X(_03797_));
 sky130_fd_sc_hd__and2_1 _16574_ (.A(_13578_),
    .B(_02422_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_1 _16575_ (.A(_13578_),
    .B(_02411_),
    .X(_03795_));
 sky130_vsdinv _16576_ (.A(\count_cycle[54] ),
    .Y(_13579_));
 sky130_fd_sc_hd__inv_2 _16577_ (.A(\count_cycle[11] ),
    .Y(_01859_));
 sky130_fd_sc_hd__inv_2 _16578_ (.A(\count_cycle[12] ),
    .Y(_01872_));
 sky130_fd_sc_hd__inv_2 _16579_ (.A(\count_cycle[7] ),
    .Y(_01806_));
 sky130_fd_sc_hd__inv_2 _16580_ (.A(\count_cycle[8] ),
    .Y(_01820_));
 sky130_fd_sc_hd__inv_2 _16581_ (.A(\count_cycle[3] ),
    .Y(_01754_));
 sky130_fd_sc_hd__inv_2 _16582_ (.A(\count_cycle[4] ),
    .Y(_01767_));
 sky130_fd_sc_hd__nand3_4 _16583_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .Y(_13580_));
 sky130_fd_sc_hd__nor3_4 _16584_ (.A(_01754_),
    .B(_01767_),
    .C(_13580_),
    .Y(_13581_));
 sky130_fd_sc_hd__nand3_4 _16585_ (.A(_13581_),
    .B(\count_cycle[5] ),
    .C(\count_cycle[6] ),
    .Y(_13582_));
 sky130_fd_sc_hd__nor3_4 _16586_ (.A(_01806_),
    .B(_01820_),
    .C(_13582_),
    .Y(_13583_));
 sky130_fd_sc_hd__nand3_4 _16587_ (.A(_13583_),
    .B(\count_cycle[9] ),
    .C(\count_cycle[10] ),
    .Y(_13584_));
 sky130_fd_sc_hd__nor3_4 _16588_ (.A(_01859_),
    .B(_01872_),
    .C(_13584_),
    .Y(_13585_));
 sky130_fd_sc_hd__and4_1 _16589_ (.A(_13585_),
    .B(\count_cycle[13] ),
    .C(\count_cycle[14] ),
    .D(\count_cycle[15] ),
    .X(_13586_));
 sky130_fd_sc_hd__and4_1 _16590_ (.A(_13586_),
    .B(\count_cycle[16] ),
    .C(\count_cycle[17] ),
    .D(\count_cycle[18] ),
    .X(_13587_));
 sky130_fd_sc_hd__clkbuf_2 _16591_ (.A(\count_cycle[19] ),
    .X(_13588_));
 sky130_fd_sc_hd__and4_1 _16592_ (.A(_13587_),
    .B(_13588_),
    .C(\count_cycle[20] ),
    .D(\count_cycle[21] ),
    .X(_13589_));
 sky130_fd_sc_hd__clkbuf_2 _16593_ (.A(\count_cycle[22] ),
    .X(_13590_));
 sky130_fd_sc_hd__and4_1 _16594_ (.A(_13589_),
    .B(_13590_),
    .C(\count_cycle[23] ),
    .D(\count_cycle[24] ),
    .X(_13591_));
 sky130_fd_sc_hd__and4_1 _16595_ (.A(_13591_),
    .B(\count_cycle[25] ),
    .C(\count_cycle[26] ),
    .D(\count_cycle[27] ),
    .X(_13592_));
 sky130_fd_sc_hd__and4_1 _16596_ (.A(_13592_),
    .B(\count_cycle[28] ),
    .C(\count_cycle[29] ),
    .D(\count_cycle[30] ),
    .X(_13593_));
 sky130_fd_sc_hd__clkbuf_2 _16597_ (.A(\count_cycle[31] ),
    .X(_13594_));
 sky130_fd_sc_hd__and4_1 _16598_ (.A(_13593_),
    .B(\count_cycle[32] ),
    .C(\count_cycle[33] ),
    .D(_13594_),
    .X(_13595_));
 sky130_fd_sc_hd__clkbuf_2 _16599_ (.A(\count_cycle[34] ),
    .X(_13596_));
 sky130_fd_sc_hd__and4_1 _16600_ (.A(_13595_),
    .B(_13596_),
    .C(\count_cycle[35] ),
    .D(\count_cycle[36] ),
    .X(_13597_));
 sky130_fd_sc_hd__and4_1 _16601_ (.A(_13597_),
    .B(\count_cycle[37] ),
    .C(\count_cycle[38] ),
    .D(\count_cycle[39] ),
    .X(_13598_));
 sky130_fd_sc_hd__clkbuf_2 _16602_ (.A(\count_cycle[40] ),
    .X(_13599_));
 sky130_fd_sc_hd__and4_1 _16603_ (.A(_13598_),
    .B(_13599_),
    .C(\count_cycle[41] ),
    .D(\count_cycle[42] ),
    .X(_13600_));
 sky130_fd_sc_hd__and4_1 _16604_ (.A(_13600_),
    .B(\count_cycle[43] ),
    .C(\count_cycle[44] ),
    .D(\count_cycle[45] ),
    .X(_13601_));
 sky130_fd_sc_hd__clkbuf_2 _16605_ (.A(\count_cycle[46] ),
    .X(_13602_));
 sky130_fd_sc_hd__and4_2 _16606_ (.A(_13601_),
    .B(_13602_),
    .C(\count_cycle[47] ),
    .D(\count_cycle[48] ),
    .X(_13603_));
 sky130_fd_sc_hd__clkbuf_2 _16607_ (.A(\count_cycle[50] ),
    .X(_13604_));
 sky130_fd_sc_hd__and4_2 _16608_ (.A(_13603_),
    .B(\count_cycle[49] ),
    .C(_13604_),
    .D(\count_cycle[51] ),
    .X(_13605_));
 sky130_fd_sc_hd__nand3_4 _16609_ (.A(_13605_),
    .B(\count_cycle[52] ),
    .C(\count_cycle[53] ),
    .Y(_13606_));
 sky130_fd_sc_hd__nor2_4 _16610_ (.A(_13579_),
    .B(_13606_),
    .Y(_13607_));
 sky130_fd_sc_hd__and4_1 _16611_ (.A(_13607_),
    .B(\count_cycle[55] ),
    .C(\count_cycle[56] ),
    .D(\count_cycle[57] ),
    .X(_13608_));
 sky130_fd_sc_hd__and4_1 _16612_ (.A(_13608_),
    .B(\count_cycle[58] ),
    .C(\count_cycle[59] ),
    .D(\count_cycle[60] ),
    .X(_13609_));
 sky130_fd_sc_hd__and4_1 _16613_ (.A(_13609_),
    .B(\count_cycle[61] ),
    .C(\count_cycle[62] ),
    .D(\count_cycle[63] ),
    .X(_13610_));
 sky130_fd_sc_hd__nor2_2 _16614_ (.A(_01859_),
    .B(_13584_),
    .Y(_13611_));
 sky130_fd_sc_hd__and4_1 _16615_ (.A(_13611_),
    .B(\count_cycle[12] ),
    .C(\count_cycle[13] ),
    .D(\count_cycle[14] ),
    .X(_13612_));
 sky130_fd_sc_hd__clkbuf_2 _16616_ (.A(\count_cycle[16] ),
    .X(_13613_));
 sky130_fd_sc_hd__and4_1 _16617_ (.A(_13612_),
    .B(\count_cycle[15] ),
    .C(_13613_),
    .D(\count_cycle[17] ),
    .X(_13614_));
 sky130_fd_sc_hd__and4_1 _16618_ (.A(_13614_),
    .B(\count_cycle[18] ),
    .C(\count_cycle[19] ),
    .D(\count_cycle[20] ),
    .X(_13615_));
 sky130_fd_sc_hd__and4_1 _16619_ (.A(_13615_),
    .B(\count_cycle[21] ),
    .C(\count_cycle[22] ),
    .D(\count_cycle[23] ),
    .X(_13616_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16620_ (.A(\count_cycle[24] ),
    .X(_13617_));
 sky130_fd_sc_hd__and4_1 _16621_ (.A(_13616_),
    .B(_13617_),
    .C(\count_cycle[25] ),
    .D(\count_cycle[26] ),
    .X(_13618_));
 sky130_fd_sc_hd__and4_1 _16622_ (.A(_13618_),
    .B(\count_cycle[27] ),
    .C(\count_cycle[28] ),
    .D(\count_cycle[29] ),
    .X(_13619_));
 sky130_fd_sc_hd__and4_1 _16623_ (.A(_13619_),
    .B(\count_cycle[32] ),
    .C(\count_cycle[30] ),
    .D(\count_cycle[31] ),
    .X(_13620_));
 sky130_fd_sc_hd__and4_1 _16624_ (.A(_13620_),
    .B(\count_cycle[33] ),
    .C(\count_cycle[34] ),
    .D(\count_cycle[35] ),
    .X(_13621_));
 sky130_fd_sc_hd__and4_1 _16625_ (.A(_13621_),
    .B(\count_cycle[36] ),
    .C(\count_cycle[37] ),
    .D(\count_cycle[38] ),
    .X(_13622_));
 sky130_fd_sc_hd__clkbuf_2 _16626_ (.A(\count_cycle[39] ),
    .X(_13623_));
 sky130_fd_sc_hd__and4_1 _16627_ (.A(_13622_),
    .B(_13623_),
    .C(\count_cycle[40] ),
    .D(\count_cycle[41] ),
    .X(_13624_));
 sky130_fd_sc_hd__and4_1 _16628_ (.A(_13624_),
    .B(\count_cycle[42] ),
    .C(\count_cycle[43] ),
    .D(\count_cycle[44] ),
    .X(_13625_));
 sky130_fd_sc_hd__clkbuf_2 _16629_ (.A(\count_cycle[45] ),
    .X(_13626_));
 sky130_fd_sc_hd__and4_1 _16630_ (.A(_13625_),
    .B(_13626_),
    .C(\count_cycle[46] ),
    .D(\count_cycle[47] ),
    .X(_13627_));
 sky130_fd_sc_hd__clkbuf_2 _16631_ (.A(\count_cycle[48] ),
    .X(_13628_));
 sky130_fd_sc_hd__and4_1 _16632_ (.A(_13627_),
    .B(_13628_),
    .C(\count_cycle[49] ),
    .D(\count_cycle[50] ),
    .X(_13629_));
 sky130_fd_sc_hd__and4_1 _16633_ (.A(_13629_),
    .B(\count_cycle[51] ),
    .C(\count_cycle[52] ),
    .D(\count_cycle[53] ),
    .X(_13630_));
 sky130_fd_sc_hd__and4_1 _16634_ (.A(_13630_),
    .B(\count_cycle[54] ),
    .C(\count_cycle[55] ),
    .D(\count_cycle[56] ),
    .X(_13631_));
 sky130_fd_sc_hd__and4_1 _16635_ (.A(_13631_),
    .B(\count_cycle[57] ),
    .C(\count_cycle[58] ),
    .D(\count_cycle[59] ),
    .X(_13632_));
 sky130_fd_sc_hd__and4_1 _16636_ (.A(_13632_),
    .B(\count_cycle[60] ),
    .C(\count_cycle[61] ),
    .D(\count_cycle[62] ),
    .X(_13633_));
 sky130_fd_sc_hd__o21bai_1 _16637_ (.A1(\count_cycle[63] ),
    .A2(_13633_),
    .B1_N(_12814_),
    .Y(_13634_));
 sky130_fd_sc_hd__nor2_1 _16638_ (.A(_13610_),
    .B(_13634_),
    .Y(_03794_));
 sky130_fd_sc_hd__clkbuf_2 _16639_ (.A(\count_cycle[59] ),
    .X(_13635_));
 sky130_fd_sc_hd__clkbuf_2 _16640_ (.A(\count_cycle[55] ),
    .X(_13636_));
 sky130_fd_sc_hd__nor3b_4 _16641_ (.A(_13579_),
    .B(_13606_),
    .C_N(_13636_),
    .Y(_13637_));
 sky130_fd_sc_hd__clkbuf_2 _16642_ (.A(\count_cycle[57] ),
    .X(_13638_));
 sky130_fd_sc_hd__and4_1 _16643_ (.A(_13637_),
    .B(\count_cycle[56] ),
    .C(_13638_),
    .D(\count_cycle[58] ),
    .X(_13639_));
 sky130_fd_sc_hd__clkbuf_2 _16644_ (.A(\count_cycle[60] ),
    .X(_13640_));
 sky130_fd_sc_hd__a41oi_1 _16645_ (.A1(_13635_),
    .A2(_13639_),
    .A3(_13640_),
    .A4(\count_cycle[61] ),
    .B1(\count_cycle[62] ),
    .Y(_13641_));
 sky130_fd_sc_hd__nor3_1 _16646_ (.A(_13452_),
    .B(_13641_),
    .C(_13633_),
    .Y(_03793_));
 sky130_fd_sc_hd__clkbuf_2 _16647_ (.A(\count_cycle[58] ),
    .X(_13642_));
 sky130_fd_sc_hd__a41oi_1 _16648_ (.A1(_13642_),
    .A2(_13608_),
    .A3(_13635_),
    .A4(_13640_),
    .B1(\count_cycle[61] ),
    .Y(_13643_));
 sky130_fd_sc_hd__and4_1 _16649_ (.A(_13639_),
    .B(_13635_),
    .C(_13640_),
    .D(\count_cycle[61] ),
    .X(_13644_));
 sky130_fd_sc_hd__nor3_1 _16650_ (.A(_13452_),
    .B(_13643_),
    .C(_13644_),
    .Y(_03792_));
 sky130_fd_sc_hd__buf_2 _16651_ (.A(_12870_),
    .X(_13645_));
 sky130_fd_sc_hd__a41oi_1 _16652_ (.A1(_13642_),
    .A2(_13608_),
    .A3(_13635_),
    .A4(_13640_),
    .B1(_13645_),
    .Y(_13646_));
 sky130_fd_sc_hd__o21a_1 _16653_ (.A1(_13640_),
    .A2(_13632_),
    .B1(_13646_),
    .X(_03791_));
 sky130_fd_sc_hd__clkbuf_2 _16654_ (.A(\count_cycle[56] ),
    .X(_13647_));
 sky130_fd_sc_hd__a41oi_2 _16655_ (.A1(_13647_),
    .A2(_13637_),
    .A3(_13638_),
    .A4(_13642_),
    .B1(_13635_),
    .Y(_13648_));
 sky130_fd_sc_hd__nor3_2 _16656_ (.A(_13452_),
    .B(_13648_),
    .C(_13632_),
    .Y(_03790_));
 sky130_fd_sc_hd__a41oi_1 _16657_ (.A1(_13647_),
    .A2(_13637_),
    .A3(_13638_),
    .A4(_13642_),
    .B1(_13645_),
    .Y(_13649_));
 sky130_fd_sc_hd__o21a_1 _16658_ (.A1(_13642_),
    .A2(_13608_),
    .B1(_13649_),
    .X(_03789_));
 sky130_fd_sc_hd__a41oi_1 _16659_ (.A1(_13636_),
    .A2(_13607_),
    .A3(_13647_),
    .A4(_13638_),
    .B1(_13645_),
    .Y(_13650_));
 sky130_fd_sc_hd__o21a_1 _16660_ (.A1(_13638_),
    .A2(_13631_),
    .B1(_13650_),
    .X(_03788_));
 sky130_fd_sc_hd__buf_2 _16661_ (.A(_12870_),
    .X(_13651_));
 sky130_fd_sc_hd__a31oi_1 _16662_ (.A1(_13607_),
    .A2(_13636_),
    .A3(_13647_),
    .B1(_13651_),
    .Y(_13652_));
 sky130_fd_sc_hd__o21a_1 _16663_ (.A1(_13647_),
    .A2(_13637_),
    .B1(_13652_),
    .X(_03787_));
 sky130_fd_sc_hd__a31oi_1 _16664_ (.A1(_13630_),
    .A2(\count_cycle[54] ),
    .A3(_13636_),
    .B1(_13651_),
    .Y(_13653_));
 sky130_fd_sc_hd__o21a_1 _16665_ (.A1(_13636_),
    .A2(_13607_),
    .B1(_13653_),
    .X(_03786_));
 sky130_fd_sc_hd__clkbuf_2 _16666_ (.A(\count_cycle[52] ),
    .X(_13654_));
 sky130_fd_sc_hd__a31oi_1 _16667_ (.A1(_13605_),
    .A2(_13654_),
    .A3(\count_cycle[53] ),
    .B1(\count_cycle[54] ),
    .Y(_13655_));
 sky130_fd_sc_hd__nor3_1 _16668_ (.A(_13452_),
    .B(_13655_),
    .C(_13607_),
    .Y(_03785_));
 sky130_fd_sc_hd__clkbuf_2 _16669_ (.A(\count_cycle[51] ),
    .X(_13656_));
 sky130_fd_sc_hd__and3_1 _16670_ (.A(_13629_),
    .B(_13656_),
    .C(_13654_),
    .X(_13657_));
 sky130_fd_sc_hd__a31oi_1 _16671_ (.A1(_13605_),
    .A2(_13654_),
    .A3(\count_cycle[53] ),
    .B1(_13651_),
    .Y(_13658_));
 sky130_fd_sc_hd__o21a_1 _16672_ (.A1(\count_cycle[53] ),
    .A2(_13657_),
    .B1(_13658_),
    .X(_03784_));
 sky130_fd_sc_hd__nand3_1 _16673_ (.A(_13629_),
    .B(_13656_),
    .C(_13654_),
    .Y(_13659_));
 sky130_fd_sc_hd__a41o_1 _16674_ (.A1(_13603_),
    .A2(\count_cycle[49] ),
    .A3(_13604_),
    .A4(_13656_),
    .B1(_13654_),
    .X(_13660_));
 sky130_fd_sc_hd__and3_1 _16675_ (.A(_13659_),
    .B(_13660_),
    .C(_13542_),
    .X(_03783_));
 sky130_fd_sc_hd__clkbuf_2 _16676_ (.A(\count_cycle[49] ),
    .X(_13661_));
 sky130_fd_sc_hd__a41oi_1 _16677_ (.A1(_13661_),
    .A2(_13603_),
    .A3(_13604_),
    .A4(_13656_),
    .B1(_13645_),
    .Y(_13662_));
 sky130_fd_sc_hd__o21a_1 _16678_ (.A1(_13656_),
    .A2(_13629_),
    .B1(_13662_),
    .X(_03782_));
 sky130_fd_sc_hd__and3_1 _16679_ (.A(_13627_),
    .B(_13628_),
    .C(_13661_),
    .X(_13663_));
 sky130_fd_sc_hd__a31oi_1 _16680_ (.A1(_13603_),
    .A2(_13661_),
    .A3(_13604_),
    .B1(_13651_),
    .Y(_13664_));
 sky130_fd_sc_hd__o21a_1 _16681_ (.A1(_13604_),
    .A2(_13663_),
    .B1(_13664_),
    .X(_03781_));
 sky130_fd_sc_hd__a31oi_1 _16682_ (.A1(_13627_),
    .A2(_13628_),
    .A3(_13661_),
    .B1(_13651_),
    .Y(_13665_));
 sky130_fd_sc_hd__o21a_1 _16683_ (.A1(_13661_),
    .A2(_13603_),
    .B1(_13665_),
    .X(_03780_));
 sky130_fd_sc_hd__a41oi_1 _16684_ (.A1(_13602_),
    .A2(_13601_),
    .A3(\count_cycle[47] ),
    .A4(_13628_),
    .B1(_13645_),
    .Y(_13666_));
 sky130_fd_sc_hd__o21a_1 _16685_ (.A1(_13628_),
    .A2(_13627_),
    .B1(_13666_),
    .X(_03779_));
 sky130_fd_sc_hd__a31oi_1 _16686_ (.A1(_13625_),
    .A2(_13626_),
    .A3(_13602_),
    .B1(\count_cycle[47] ),
    .Y(_13667_));
 sky130_fd_sc_hd__nor3_1 _16687_ (.A(_13452_),
    .B(_13667_),
    .C(_13627_),
    .Y(_03778_));
 sky130_fd_sc_hd__a31oi_1 _16688_ (.A1(_13625_),
    .A2(_13626_),
    .A3(_13602_),
    .B1(_13651_),
    .Y(_13668_));
 sky130_fd_sc_hd__o21a_1 _16689_ (.A1(_13602_),
    .A2(_13601_),
    .B1(_13668_),
    .X(_03777_));
 sky130_fd_sc_hd__clkbuf_2 _16690_ (.A(\count_cycle[43] ),
    .X(_13669_));
 sky130_fd_sc_hd__a41oi_1 _16691_ (.A1(_13669_),
    .A2(_13600_),
    .A3(\count_cycle[44] ),
    .A4(_13626_),
    .B1(_12871_),
    .Y(_13670_));
 sky130_fd_sc_hd__o21a_1 _16692_ (.A1(_13626_),
    .A2(_13625_),
    .B1(_13670_),
    .X(_03776_));
 sky130_fd_sc_hd__and3_1 _16693_ (.A(_13624_),
    .B(\count_cycle[42] ),
    .C(_13669_),
    .X(_13671_));
 sky130_fd_sc_hd__buf_2 _16694_ (.A(_12870_),
    .X(_13672_));
 sky130_fd_sc_hd__a31oi_1 _16695_ (.A1(_13600_),
    .A2(_13669_),
    .A3(\count_cycle[44] ),
    .B1(_13672_),
    .Y(_13673_));
 sky130_fd_sc_hd__o21a_1 _16696_ (.A1(\count_cycle[44] ),
    .A2(_13671_),
    .B1(_13673_),
    .X(_03775_));
 sky130_fd_sc_hd__a31oi_1 _16697_ (.A1(_13624_),
    .A2(\count_cycle[42] ),
    .A3(_13669_),
    .B1(_13672_),
    .Y(_13674_));
 sky130_fd_sc_hd__o21a_1 _16698_ (.A1(_13669_),
    .A2(_13600_),
    .B1(_13674_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_2 _16699_ (.A(_13321_),
    .X(_13675_));
 sky130_fd_sc_hd__a31oi_1 _16700_ (.A1(_13598_),
    .A2(_13599_),
    .A3(\count_cycle[41] ),
    .B1(\count_cycle[42] ),
    .Y(_13676_));
 sky130_fd_sc_hd__nor3_1 _16701_ (.A(_13675_),
    .B(_13676_),
    .C(_13600_),
    .Y(_03773_));
 sky130_fd_sc_hd__a31oi_1 _16702_ (.A1(_13622_),
    .A2(_13623_),
    .A3(_13599_),
    .B1(\count_cycle[41] ),
    .Y(_13677_));
 sky130_fd_sc_hd__nor3_1 _16703_ (.A(_13675_),
    .B(_13677_),
    .C(_13624_),
    .Y(_03772_));
 sky130_fd_sc_hd__nand3_1 _16704_ (.A(_13622_),
    .B(_13623_),
    .C(_13599_),
    .Y(_13678_));
 sky130_fd_sc_hd__clkbuf_2 _16705_ (.A(\count_cycle[37] ),
    .X(_13679_));
 sky130_fd_sc_hd__a41o_1 _16706_ (.A1(_13597_),
    .A2(_13679_),
    .A3(\count_cycle[38] ),
    .A4(_13623_),
    .B1(_13599_),
    .X(_13680_));
 sky130_fd_sc_hd__and3_1 _16707_ (.A(_13678_),
    .B(_13680_),
    .C(_13542_),
    .X(_03771_));
 sky130_fd_sc_hd__a31oi_1 _16708_ (.A1(_13597_),
    .A2(_13679_),
    .A3(\count_cycle[38] ),
    .B1(_13623_),
    .Y(_13681_));
 sky130_fd_sc_hd__nor3_1 _16709_ (.A(_13675_),
    .B(_13681_),
    .C(_13598_),
    .Y(_03770_));
 sky130_fd_sc_hd__a31oi_1 _16710_ (.A1(_13621_),
    .A2(\count_cycle[36] ),
    .A3(_13679_),
    .B1(\count_cycle[38] ),
    .Y(_13682_));
 sky130_fd_sc_hd__nor3_1 _16711_ (.A(_13675_),
    .B(_13682_),
    .C(_13622_),
    .Y(_03769_));
 sky130_fd_sc_hd__a31oi_1 _16712_ (.A1(_13621_),
    .A2(\count_cycle[36] ),
    .A3(_13679_),
    .B1(_13672_),
    .Y(_13683_));
 sky130_fd_sc_hd__o21a_1 _16713_ (.A1(_13679_),
    .A2(_13597_),
    .B1(_13683_),
    .X(_03768_));
 sky130_fd_sc_hd__a31oi_1 _16714_ (.A1(_13595_),
    .A2(_13596_),
    .A3(\count_cycle[35] ),
    .B1(\count_cycle[36] ),
    .Y(_13684_));
 sky130_fd_sc_hd__nor3_1 _16715_ (.A(_13675_),
    .B(_13684_),
    .C(_13597_),
    .Y(_03767_));
 sky130_fd_sc_hd__a31oi_1 _16716_ (.A1(_13620_),
    .A2(\count_cycle[33] ),
    .A3(_13596_),
    .B1(\count_cycle[35] ),
    .Y(_13685_));
 sky130_fd_sc_hd__nor3_1 _16717_ (.A(_13675_),
    .B(_13685_),
    .C(_13621_),
    .Y(_03766_));
 sky130_fd_sc_hd__a31oi_1 _16718_ (.A1(_13620_),
    .A2(\count_cycle[33] ),
    .A3(_13596_),
    .B1(_13672_),
    .Y(_13686_));
 sky130_fd_sc_hd__o21a_1 _16719_ (.A1(_13596_),
    .A2(_13595_),
    .B1(_13686_),
    .X(_03765_));
 sky130_fd_sc_hd__buf_2 _16720_ (.A(_13321_),
    .X(_13687_));
 sky130_fd_sc_hd__a31oi_1 _16721_ (.A1(_13593_),
    .A2(\count_cycle[32] ),
    .A3(_13594_),
    .B1(\count_cycle[33] ),
    .Y(_13688_));
 sky130_fd_sc_hd__nor3_1 _16722_ (.A(_13687_),
    .B(_13688_),
    .C(_13595_),
    .Y(_03764_));
 sky130_fd_sc_hd__a31oi_1 _16723_ (.A1(_13619_),
    .A2(\count_cycle[30] ),
    .A3(_13594_),
    .B1(\count_cycle[32] ),
    .Y(_13689_));
 sky130_fd_sc_hd__nor3_1 _16724_ (.A(_13687_),
    .B(_13689_),
    .C(_13620_),
    .Y(_03763_));
 sky130_fd_sc_hd__a31oi_1 _16725_ (.A1(_13619_),
    .A2(\count_cycle[30] ),
    .A3(_13594_),
    .B1(_13672_),
    .Y(_13690_));
 sky130_fd_sc_hd__o21a_1 _16726_ (.A1(_13594_),
    .A2(_13593_),
    .B1(_13690_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_2 _16727_ (.A(\count_cycle[28] ),
    .X(_13691_));
 sky130_fd_sc_hd__a31oi_1 _16728_ (.A1(_13592_),
    .A2(_13691_),
    .A3(\count_cycle[29] ),
    .B1(\count_cycle[30] ),
    .Y(_13692_));
 sky130_fd_sc_hd__nor3_1 _16729_ (.A(_13687_),
    .B(_13692_),
    .C(_13593_),
    .Y(_03761_));
 sky130_fd_sc_hd__and3_1 _16730_ (.A(_13618_),
    .B(\count_cycle[27] ),
    .C(_13691_),
    .X(_13693_));
 sky130_fd_sc_hd__a31oi_1 _16731_ (.A1(_13592_),
    .A2(_13691_),
    .A3(\count_cycle[29] ),
    .B1(_13672_),
    .Y(_13694_));
 sky130_fd_sc_hd__o21a_1 _16732_ (.A1(\count_cycle[29] ),
    .A2(_13693_),
    .B1(_13694_),
    .X(_03760_));
 sky130_fd_sc_hd__buf_2 _16733_ (.A(_12870_),
    .X(_13695_));
 sky130_fd_sc_hd__a31oi_1 _16734_ (.A1(_13618_),
    .A2(\count_cycle[27] ),
    .A3(_13691_),
    .B1(_13695_),
    .Y(_13696_));
 sky130_fd_sc_hd__o21a_1 _16735_ (.A1(_13691_),
    .A2(_13592_),
    .B1(_13696_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_2 _16736_ (.A(\count_cycle[25] ),
    .X(_13697_));
 sky130_fd_sc_hd__a31oi_1 _16737_ (.A1(_13591_),
    .A2(_13697_),
    .A3(\count_cycle[26] ),
    .B1(\count_cycle[27] ),
    .Y(_13698_));
 sky130_fd_sc_hd__nor3_1 _16738_ (.A(_13687_),
    .B(_13698_),
    .C(_13592_),
    .Y(_03758_));
 sky130_fd_sc_hd__and3_1 _16739_ (.A(_13616_),
    .B(_13617_),
    .C(_13697_),
    .X(_13699_));
 sky130_fd_sc_hd__a31oi_1 _16740_ (.A1(_13591_),
    .A2(_13697_),
    .A3(\count_cycle[26] ),
    .B1(_13695_),
    .Y(_13700_));
 sky130_fd_sc_hd__o21a_1 _16741_ (.A1(\count_cycle[26] ),
    .A2(_13699_),
    .B1(_13700_),
    .X(_03757_));
 sky130_fd_sc_hd__a31oi_1 _16742_ (.A1(_13616_),
    .A2(_13617_),
    .A3(_13697_),
    .B1(_13695_),
    .Y(_13701_));
 sky130_fd_sc_hd__o21a_1 _16743_ (.A1(_13697_),
    .A2(_13591_),
    .B1(_13701_),
    .X(_03756_));
 sky130_fd_sc_hd__a41oi_1 _16744_ (.A1(_13590_),
    .A2(_13589_),
    .A3(\count_cycle[23] ),
    .A4(_13617_),
    .B1(_12871_),
    .Y(_13702_));
 sky130_fd_sc_hd__o21a_1 _16745_ (.A1(_13617_),
    .A2(_13616_),
    .B1(_13702_),
    .X(_03755_));
 sky130_fd_sc_hd__a31oi_1 _16746_ (.A1(_13615_),
    .A2(\count_cycle[21] ),
    .A3(_13590_),
    .B1(\count_cycle[23] ),
    .Y(_13703_));
 sky130_fd_sc_hd__nor3_1 _16747_ (.A(_13687_),
    .B(_13703_),
    .C(_13616_),
    .Y(_03754_));
 sky130_fd_sc_hd__a31oi_1 _16748_ (.A1(_13615_),
    .A2(\count_cycle[21] ),
    .A3(_13590_),
    .B1(_13695_),
    .Y(_13704_));
 sky130_fd_sc_hd__o21a_1 _16749_ (.A1(_13590_),
    .A2(_13589_),
    .B1(_13704_),
    .X(_03753_));
 sky130_fd_sc_hd__a31oi_1 _16750_ (.A1(_13587_),
    .A2(_13588_),
    .A3(\count_cycle[20] ),
    .B1(\count_cycle[21] ),
    .Y(_13705_));
 sky130_fd_sc_hd__nor3_1 _16751_ (.A(_13687_),
    .B(_13705_),
    .C(_13589_),
    .Y(_03752_));
 sky130_fd_sc_hd__buf_2 _16752_ (.A(_13321_),
    .X(_13706_));
 sky130_fd_sc_hd__a31oi_1 _16753_ (.A1(_13614_),
    .A2(\count_cycle[18] ),
    .A3(_13588_),
    .B1(\count_cycle[20] ),
    .Y(_13707_));
 sky130_fd_sc_hd__nor3_1 _16754_ (.A(_13706_),
    .B(_13707_),
    .C(_13615_),
    .Y(_03751_));
 sky130_fd_sc_hd__a31oi_1 _16755_ (.A1(_13614_),
    .A2(\count_cycle[18] ),
    .A3(_13588_),
    .B1(_13695_),
    .Y(_13708_));
 sky130_fd_sc_hd__o21a_1 _16756_ (.A1(_13588_),
    .A2(_13587_),
    .B1(_13708_),
    .X(_03750_));
 sky130_fd_sc_hd__a31oi_1 _16757_ (.A1(_13586_),
    .A2(_13613_),
    .A3(\count_cycle[17] ),
    .B1(\count_cycle[18] ),
    .Y(_13709_));
 sky130_fd_sc_hd__nor3_1 _16758_ (.A(_13706_),
    .B(_13709_),
    .C(_13587_),
    .Y(_03749_));
 sky130_fd_sc_hd__a31oi_1 _16759_ (.A1(_13612_),
    .A2(\count_cycle[15] ),
    .A3(_13613_),
    .B1(\count_cycle[17] ),
    .Y(_13710_));
 sky130_fd_sc_hd__nor3_1 _16760_ (.A(_13706_),
    .B(_13710_),
    .C(_13614_),
    .Y(_03748_));
 sky130_fd_sc_hd__a31oi_1 _16761_ (.A1(_13612_),
    .A2(\count_cycle[15] ),
    .A3(_13613_),
    .B1(_13695_),
    .Y(_13711_));
 sky130_fd_sc_hd__o21a_1 _16762_ (.A1(_13613_),
    .A2(_13586_),
    .B1(_13711_),
    .X(_03747_));
 sky130_fd_sc_hd__a31oi_1 _16763_ (.A1(_13585_),
    .A2(\count_cycle[13] ),
    .A3(\count_cycle[14] ),
    .B1(\count_cycle[15] ),
    .Y(_13712_));
 sky130_fd_sc_hd__nor3_1 _16764_ (.A(_13706_),
    .B(_13712_),
    .C(_13586_),
    .Y(_03746_));
 sky130_fd_sc_hd__a31oi_1 _16765_ (.A1(_13611_),
    .A2(\count_cycle[12] ),
    .A3(\count_cycle[13] ),
    .B1(\count_cycle[14] ),
    .Y(_13713_));
 sky130_fd_sc_hd__nor3_1 _16766_ (.A(_13706_),
    .B(_13713_),
    .C(_13612_),
    .Y(_03745_));
 sky130_fd_sc_hd__inv_2 _16767_ (.A(\count_cycle[13] ),
    .Y(_01885_));
 sky130_vsdinv _16768_ (.A(_13585_),
    .Y(_13714_));
 sky130_fd_sc_hd__o41ai_1 _16769_ (.A1(_01859_),
    .A2(_01872_),
    .A3(_01885_),
    .A4(_13584_),
    .B1(_13333_),
    .Y(_13715_));
 sky130_fd_sc_hd__a21oi_1 _16770_ (.A1(_01885_),
    .A2(_13714_),
    .B1(_13715_),
    .Y(_03744_));
 sky130_fd_sc_hd__a41oi_1 _16771_ (.A1(\count_cycle[9] ),
    .A2(_13583_),
    .A3(\count_cycle[10] ),
    .A4(\count_cycle[11] ),
    .B1(\count_cycle[12] ),
    .Y(_13716_));
 sky130_fd_sc_hd__nor3_1 _16772_ (.A(_13706_),
    .B(_13716_),
    .C(_13585_),
    .Y(_03743_));
 sky130_fd_sc_hd__buf_4 _16773_ (.A(_12814_),
    .X(_13717_));
 sky130_fd_sc_hd__a31oi_1 _16774_ (.A1(_13583_),
    .A2(\count_cycle[9] ),
    .A3(\count_cycle[10] ),
    .B1(\count_cycle[11] ),
    .Y(_13718_));
 sky130_fd_sc_hd__nor3_1 _16775_ (.A(_13717_),
    .B(_13718_),
    .C(_13611_),
    .Y(_03742_));
 sky130_fd_sc_hd__inv_2 _16776_ (.A(\count_cycle[9] ),
    .Y(_01833_));
 sky130_fd_sc_hd__inv_2 _16777_ (.A(\count_cycle[10] ),
    .Y(_01846_));
 sky130_fd_sc_hd__o41ai_1 _16778_ (.A1(_01806_),
    .A2(_01820_),
    .A3(_01833_),
    .A4(_13582_),
    .B1(_01846_),
    .Y(_13719_));
 sky130_fd_sc_hd__and3_1 _16779_ (.A(_13719_),
    .B(_13584_),
    .C(_13329_),
    .X(_03741_));
 sky130_fd_sc_hd__inv_2 _16780_ (.A(\count_cycle[6] ),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_2 _16781_ (.A(_01754_),
    .B(_13580_),
    .Y(_13720_));
 sky130_fd_sc_hd__nand3_4 _16782_ (.A(_13720_),
    .B(\count_cycle[4] ),
    .C(\count_cycle[5] ),
    .Y(_13721_));
 sky130_fd_sc_hd__nor3_4 _16783_ (.A(_01793_),
    .B(_01806_),
    .C(_13721_),
    .Y(_13722_));
 sky130_fd_sc_hd__a31oi_1 _16784_ (.A1(_13722_),
    .A2(\count_cycle[8] ),
    .A3(\count_cycle[9] ),
    .B1(_13645_),
    .Y(_13723_));
 sky130_fd_sc_hd__o21a_1 _16785_ (.A1(\count_cycle[9] ),
    .A2(_13583_),
    .B1(_13723_),
    .X(_03740_));
 sky130_fd_sc_hd__a41oi_1 _16786_ (.A1(\count_cycle[5] ),
    .A2(_13581_),
    .A3(\count_cycle[6] ),
    .A4(\count_cycle[7] ),
    .B1(\count_cycle[8] ),
    .Y(_13724_));
 sky130_fd_sc_hd__nor3_1 _16787_ (.A(_13717_),
    .B(_13724_),
    .C(_13583_),
    .Y(_03739_));
 sky130_fd_sc_hd__a31oi_1 _16788_ (.A1(_13581_),
    .A2(\count_cycle[5] ),
    .A3(\count_cycle[6] ),
    .B1(\count_cycle[7] ),
    .Y(_13725_));
 sky130_fd_sc_hd__nor3_1 _16789_ (.A(_13717_),
    .B(_13725_),
    .C(_13722_),
    .Y(_03738_));
 sky130_fd_sc_hd__nand2_1 _16790_ (.A(_13582_),
    .B(_13329_),
    .Y(_13726_));
 sky130_fd_sc_hd__a21oi_1 _16791_ (.A1(_01793_),
    .A2(_13721_),
    .B1(_13726_),
    .Y(_03737_));
 sky130_fd_sc_hd__inv_2 _16792_ (.A(\count_cycle[5] ),
    .Y(_01780_));
 sky130_fd_sc_hd__o31ai_1 _16793_ (.A1(_01754_),
    .A2(_01767_),
    .A3(_13580_),
    .B1(_01780_),
    .Y(_13727_));
 sky130_fd_sc_hd__and3_1 _16794_ (.A(_13727_),
    .B(_13329_),
    .C(_13721_),
    .X(_03736_));
 sky130_fd_sc_hd__clkbuf_2 _16795_ (.A(\count_cycle[0] ),
    .X(_13728_));
 sky130_fd_sc_hd__a41oi_1 _16796_ (.A1(_13728_),
    .A2(\count_cycle[1] ),
    .A3(\count_cycle[2] ),
    .A4(\count_cycle[3] ),
    .B1(\count_cycle[4] ),
    .Y(_13729_));
 sky130_fd_sc_hd__nor3_1 _16797_ (.A(_13717_),
    .B(_13581_),
    .C(_13729_),
    .Y(_03735_));
 sky130_fd_sc_hd__a31oi_1 _16798_ (.A1(_13728_),
    .A2(\count_cycle[1] ),
    .A3(\count_cycle[2] ),
    .B1(\count_cycle[3] ),
    .Y(_13730_));
 sky130_fd_sc_hd__nor3_1 _16799_ (.A(_13717_),
    .B(_13720_),
    .C(_13730_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _16800_ (.A(_13728_),
    .B(\count_cycle[1] ),
    .Y(_13731_));
 sky130_fd_sc_hd__inv_2 _16801_ (.A(\count_cycle[2] ),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_1 _16802_ (.A(_13731_),
    .B(_01741_),
    .Y(_13732_));
 sky130_fd_sc_hd__and3_1 _16803_ (.A(_13732_),
    .B(_13329_),
    .C(_13580_),
    .X(_03733_));
 sky130_fd_sc_hd__nor2_1 _16804_ (.A(_13728_),
    .B(\count_cycle[1] ),
    .Y(_13733_));
 sky130_fd_sc_hd__nor3b_1 _16805_ (.A(_12815_),
    .B(_13733_),
    .C_N(_13731_),
    .Y(_03732_));
 sky130_vsdinv _16806_ (.A(_13728_),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2b_1 _16807_ (.A(_13728_),
    .B_N(_12650_),
    .Y(_03731_));
 sky130_fd_sc_hd__and2_1 _16808_ (.A(_13578_),
    .B(\cpu_state[0] ),
    .X(_03730_));
 sky130_fd_sc_hd__and2_1 _16809_ (.A(_13578_),
    .B(\pcpi_mul.active[0] ),
    .X(_03729_));
 sky130_fd_sc_hd__buf_1 _16810_ (.A(\cpuregs_wrdata[31] ),
    .X(_13734_));
 sky130_vsdinv _16811_ (.A(latched_branch),
    .Y(_13735_));
 sky130_vsdinv _16812_ (.A(latched_store),
    .Y(_13736_));
 sky130_fd_sc_hd__and3_1 _16813_ (.A(_12698_),
    .B(_13735_),
    .C(_13736_),
    .X(_13737_));
 sky130_fd_sc_hd__nor3_4 _16814_ (.A(\latched_rd[4] ),
    .B(\latched_rd[2] ),
    .C(\latched_rd[3] ),
    .Y(_13738_));
 sky130_fd_sc_hd__nor2_8 _16815_ (.A(\latched_rd[0] ),
    .B(\latched_rd[1] ),
    .Y(_13739_));
 sky130_fd_sc_hd__and2_2 _16816_ (.A(_13738_),
    .B(_13739_),
    .X(_13740_));
 sky130_fd_sc_hd__or4_4 _16817_ (.A(_12641_),
    .B(_12847_),
    .C(_13737_),
    .D(_13740_),
    .X(_13741_));
 sky130_fd_sc_hd__buf_2 _16818_ (.A(_13741_),
    .X(_13742_));
 sky130_fd_sc_hd__nor3b_4 _16819_ (.A(\latched_rd[0] ),
    .B(_13742_),
    .C_N(\latched_rd[1] ),
    .Y(_13743_));
 sky130_fd_sc_hd__clkbuf_4 _16820_ (.A(\latched_rd[3] ),
    .X(_13744_));
 sky130_fd_sc_hd__clkbuf_4 _16821_ (.A(\latched_rd[2] ),
    .X(_13745_));
 sky130_fd_sc_hd__nor3b_4 _16822_ (.A(\latched_rd[4] ),
    .B(_13744_),
    .C_N(_13745_),
    .Y(_13746_));
 sky130_fd_sc_hd__nand2_1 _16823_ (.A(_13743_),
    .B(_13746_),
    .Y(_13747_));
 sky130_fd_sc_hd__clkbuf_8 _16824_ (.A(_13747_),
    .X(_13748_));
 sky130_fd_sc_hd__buf_4 _16825_ (.A(_13748_),
    .X(_13749_));
 sky130_fd_sc_hd__mux2_1 _16826_ (.A0(_13734_),
    .A1(\cpuregs[6][31] ),
    .S(_13749_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_2 _16827_ (.A(\cpuregs_wrdata[30] ),
    .X(_13750_));
 sky130_fd_sc_hd__mux2_1 _16828_ (.A0(_13750_),
    .A1(\cpuregs[6][30] ),
    .S(_13749_),
    .X(_03726_));
 sky130_fd_sc_hd__clkbuf_2 _16829_ (.A(\cpuregs_wrdata[29] ),
    .X(_13751_));
 sky130_fd_sc_hd__mux2_1 _16830_ (.A0(_13751_),
    .A1(\cpuregs[6][29] ),
    .S(_13749_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_2 _16831_ (.A(\cpuregs_wrdata[28] ),
    .X(_13752_));
 sky130_fd_sc_hd__mux2_1 _16832_ (.A0(_13752_),
    .A1(\cpuregs[6][28] ),
    .S(_13749_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_2 _16833_ (.A(\cpuregs_wrdata[27] ),
    .X(_13753_));
 sky130_fd_sc_hd__mux2_1 _16834_ (.A0(_13753_),
    .A1(\cpuregs[6][27] ),
    .S(_13749_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_2 _16835_ (.A(\cpuregs_wrdata[26] ),
    .X(_13754_));
 sky130_fd_sc_hd__mux2_1 _16836_ (.A0(_13754_),
    .A1(\cpuregs[6][26] ),
    .S(_13749_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_2 _16837_ (.A(\cpuregs_wrdata[25] ),
    .X(_13755_));
 sky130_fd_sc_hd__clkbuf_4 _16838_ (.A(_13748_),
    .X(_13756_));
 sky130_fd_sc_hd__mux2_1 _16839_ (.A0(_13755_),
    .A1(\cpuregs[6][25] ),
    .S(_13756_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_2 _16840_ (.A(\cpuregs_wrdata[24] ),
    .X(_13757_));
 sky130_fd_sc_hd__mux2_1 _16841_ (.A0(_13757_),
    .A1(\cpuregs[6][24] ),
    .S(_13756_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_2 _16842_ (.A(\cpuregs_wrdata[23] ),
    .X(_13758_));
 sky130_fd_sc_hd__mux2_1 _16843_ (.A0(_13758_),
    .A1(\cpuregs[6][23] ),
    .S(_13756_),
    .X(_03719_));
 sky130_fd_sc_hd__clkbuf_2 _16844_ (.A(\cpuregs_wrdata[22] ),
    .X(_13759_));
 sky130_fd_sc_hd__mux2_1 _16845_ (.A0(_13759_),
    .A1(\cpuregs[6][22] ),
    .S(_13756_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_2 _16846_ (.A(\cpuregs_wrdata[21] ),
    .X(_13760_));
 sky130_fd_sc_hd__mux2_1 _16847_ (.A0(_13760_),
    .A1(\cpuregs[6][21] ),
    .S(_13756_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_2 _16848_ (.A(\cpuregs_wrdata[20] ),
    .X(_13761_));
 sky130_fd_sc_hd__mux2_1 _16849_ (.A0(_13761_),
    .A1(\cpuregs[6][20] ),
    .S(_13756_),
    .X(_03716_));
 sky130_fd_sc_hd__clkbuf_2 _16850_ (.A(\cpuregs_wrdata[19] ),
    .X(_13762_));
 sky130_fd_sc_hd__buf_2 _16851_ (.A(_13748_),
    .X(_13763_));
 sky130_fd_sc_hd__mux2_1 _16852_ (.A0(_13762_),
    .A1(\cpuregs[6][19] ),
    .S(_13763_),
    .X(_03715_));
 sky130_fd_sc_hd__buf_2 _16853_ (.A(\cpuregs_wrdata[18] ),
    .X(_13764_));
 sky130_fd_sc_hd__mux2_1 _16854_ (.A0(_13764_),
    .A1(\cpuregs[6][18] ),
    .S(_13763_),
    .X(_03714_));
 sky130_fd_sc_hd__buf_2 _16855_ (.A(\cpuregs_wrdata[17] ),
    .X(_13765_));
 sky130_fd_sc_hd__mux2_1 _16856_ (.A0(_13765_),
    .A1(\cpuregs[6][17] ),
    .S(_13763_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_2 _16857_ (.A(\cpuregs_wrdata[16] ),
    .X(_13766_));
 sky130_fd_sc_hd__mux2_1 _16858_ (.A0(_13766_),
    .A1(\cpuregs[6][16] ),
    .S(_13763_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_2 _16859_ (.A(\cpuregs_wrdata[15] ),
    .X(_13767_));
 sky130_fd_sc_hd__mux2_1 _16860_ (.A0(_13767_),
    .A1(\cpuregs[6][15] ),
    .S(_13763_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_2 _16861_ (.A(\cpuregs_wrdata[14] ),
    .X(_13768_));
 sky130_fd_sc_hd__mux2_1 _16862_ (.A0(_13768_),
    .A1(\cpuregs[6][14] ),
    .S(_13763_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_2 _16863_ (.A(\cpuregs_wrdata[13] ),
    .X(_13769_));
 sky130_fd_sc_hd__buf_4 _16864_ (.A(_13748_),
    .X(_13770_));
 sky130_fd_sc_hd__mux2_1 _16865_ (.A0(_13769_),
    .A1(\cpuregs[6][13] ),
    .S(_13770_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_2 _16866_ (.A(\cpuregs_wrdata[12] ),
    .X(_13771_));
 sky130_fd_sc_hd__mux2_1 _16867_ (.A0(_13771_),
    .A1(\cpuregs[6][12] ),
    .S(_13770_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_2 _16868_ (.A(\cpuregs_wrdata[11] ),
    .X(_13772_));
 sky130_fd_sc_hd__mux2_1 _16869_ (.A0(_13772_),
    .A1(\cpuregs[6][11] ),
    .S(_13770_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_2 _16870_ (.A(\cpuregs_wrdata[10] ),
    .X(_13773_));
 sky130_fd_sc_hd__mux2_1 _16871_ (.A0(_13773_),
    .A1(\cpuregs[6][10] ),
    .S(_13770_),
    .X(_03706_));
 sky130_fd_sc_hd__clkbuf_2 _16872_ (.A(\cpuregs_wrdata[9] ),
    .X(_13774_));
 sky130_fd_sc_hd__mux2_1 _16873_ (.A0(_13774_),
    .A1(\cpuregs[6][9] ),
    .S(_13770_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_2 _16874_ (.A(\cpuregs_wrdata[8] ),
    .X(_13775_));
 sky130_fd_sc_hd__mux2_1 _16875_ (.A0(_13775_),
    .A1(\cpuregs[6][8] ),
    .S(_13770_),
    .X(_03704_));
 sky130_fd_sc_hd__clkbuf_2 _16876_ (.A(\cpuregs_wrdata[7] ),
    .X(_13776_));
 sky130_fd_sc_hd__clkbuf_4 _16877_ (.A(_13747_),
    .X(_13777_));
 sky130_fd_sc_hd__mux2_1 _16878_ (.A0(_13776_),
    .A1(\cpuregs[6][7] ),
    .S(_13777_),
    .X(_03703_));
 sky130_fd_sc_hd__clkbuf_2 _16879_ (.A(\cpuregs_wrdata[6] ),
    .X(_13778_));
 sky130_fd_sc_hd__mux2_1 _16880_ (.A0(_13778_),
    .A1(\cpuregs[6][6] ),
    .S(_13777_),
    .X(_03702_));
 sky130_fd_sc_hd__clkbuf_2 _16881_ (.A(\cpuregs_wrdata[5] ),
    .X(_13779_));
 sky130_fd_sc_hd__mux2_1 _16882_ (.A0(_13779_),
    .A1(\cpuregs[6][5] ),
    .S(_13777_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_2 _16883_ (.A(\cpuregs_wrdata[4] ),
    .X(_13780_));
 sky130_fd_sc_hd__mux2_1 _16884_ (.A0(_13780_),
    .A1(\cpuregs[6][4] ),
    .S(_13777_),
    .X(_03700_));
 sky130_fd_sc_hd__clkbuf_2 _16885_ (.A(\cpuregs_wrdata[3] ),
    .X(_13781_));
 sky130_fd_sc_hd__mux2_1 _16886_ (.A0(_13781_),
    .A1(\cpuregs[6][3] ),
    .S(_13777_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_2 _16887_ (.A(\cpuregs_wrdata[2] ),
    .X(_13782_));
 sky130_fd_sc_hd__mux2_1 _16888_ (.A0(_13782_),
    .A1(\cpuregs[6][2] ),
    .S(_13777_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_2 _16889_ (.A(\cpuregs_wrdata[1] ),
    .X(_13783_));
 sky130_fd_sc_hd__mux2_1 _16890_ (.A0(_13783_),
    .A1(\cpuregs[6][1] ),
    .S(_13748_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_2 _16891_ (.A(\cpuregs_wrdata[0] ),
    .X(_13784_));
 sky130_fd_sc_hd__mux2_1 _16892_ (.A0(_13784_),
    .A1(\cpuregs[6][0] ),
    .S(_13748_),
    .X(_03696_));
 sky130_vsdinv _16893_ (.A(\latched_rd[0] ),
    .Y(_13785_));
 sky130_fd_sc_hd__nor3_4 _16894_ (.A(_13785_),
    .B(\latched_rd[1] ),
    .C(_13741_),
    .Y(_13786_));
 sky130_fd_sc_hd__nor3b_4 _16895_ (.A(\latched_rd[4] ),
    .B(_13745_),
    .C_N(_13744_),
    .Y(_13787_));
 sky130_fd_sc_hd__nand2_1 _16896_ (.A(_13786_),
    .B(_13787_),
    .Y(_13788_));
 sky130_fd_sc_hd__buf_6 _16897_ (.A(_13788_),
    .X(_13789_));
 sky130_fd_sc_hd__clkbuf_4 _16898_ (.A(_13789_),
    .X(_13790_));
 sky130_fd_sc_hd__mux2_1 _16899_ (.A0(_13734_),
    .A1(\cpuregs[9][31] ),
    .S(_13790_),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_1 _16900_ (.A0(_13750_),
    .A1(\cpuregs[9][30] ),
    .S(_13790_),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_1 _16901_ (.A0(_13751_),
    .A1(\cpuregs[9][29] ),
    .S(_13790_),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _16902_ (.A0(_13752_),
    .A1(\cpuregs[9][28] ),
    .S(_13790_),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_1 _16903_ (.A0(_13753_),
    .A1(\cpuregs[9][27] ),
    .S(_13790_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _16904_ (.A0(_13754_),
    .A1(\cpuregs[9][26] ),
    .S(_13790_),
    .X(_03690_));
 sky130_fd_sc_hd__buf_2 _16905_ (.A(_13789_),
    .X(_13791_));
 sky130_fd_sc_hd__mux2_1 _16906_ (.A0(_13755_),
    .A1(\cpuregs[9][25] ),
    .S(_13791_),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_1 _16907_ (.A0(_13757_),
    .A1(\cpuregs[9][24] ),
    .S(_13791_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _16908_ (.A0(_13758_),
    .A1(\cpuregs[9][23] ),
    .S(_13791_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _16909_ (.A0(_13759_),
    .A1(\cpuregs[9][22] ),
    .S(_13791_),
    .X(_03686_));
 sky130_fd_sc_hd__mux2_1 _16910_ (.A0(_13760_),
    .A1(\cpuregs[9][21] ),
    .S(_13791_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _16911_ (.A0(_13761_),
    .A1(\cpuregs[9][20] ),
    .S(_13791_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_4 _16912_ (.A(_13789_),
    .X(_13792_));
 sky130_fd_sc_hd__mux2_1 _16913_ (.A0(_13762_),
    .A1(\cpuregs[9][19] ),
    .S(_13792_),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_1 _16914_ (.A0(_13764_),
    .A1(\cpuregs[9][18] ),
    .S(_13792_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _16915_ (.A0(_13765_),
    .A1(\cpuregs[9][17] ),
    .S(_13792_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_1 _16916_ (.A0(_13766_),
    .A1(\cpuregs[9][16] ),
    .S(_13792_),
    .X(_03680_));
 sky130_fd_sc_hd__mux2_1 _16917_ (.A0(_13767_),
    .A1(\cpuregs[9][15] ),
    .S(_13792_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _16918_ (.A0(_13768_),
    .A1(\cpuregs[9][14] ),
    .S(_13792_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_4 _16919_ (.A(_13789_),
    .X(_13793_));
 sky130_fd_sc_hd__mux2_1 _16920_ (.A0(_13769_),
    .A1(\cpuregs[9][13] ),
    .S(_13793_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _16921_ (.A0(_13771_),
    .A1(\cpuregs[9][12] ),
    .S(_13793_),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_1 _16922_ (.A0(_13772_),
    .A1(\cpuregs[9][11] ),
    .S(_13793_),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_1 _16923_ (.A0(_13773_),
    .A1(\cpuregs[9][10] ),
    .S(_13793_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _16924_ (.A0(_13774_),
    .A1(\cpuregs[9][9] ),
    .S(_13793_),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_1 _16925_ (.A0(_13775_),
    .A1(\cpuregs[9][8] ),
    .S(_13793_),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_4 _16926_ (.A(_13788_),
    .X(_13794_));
 sky130_fd_sc_hd__mux2_1 _16927_ (.A0(_13776_),
    .A1(\cpuregs[9][7] ),
    .S(_13794_),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _16928_ (.A0(_13778_),
    .A1(\cpuregs[9][6] ),
    .S(_13794_),
    .X(_03670_));
 sky130_fd_sc_hd__mux2_1 _16929_ (.A0(_13779_),
    .A1(\cpuregs[9][5] ),
    .S(_13794_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _16930_ (.A0(_13780_),
    .A1(\cpuregs[9][4] ),
    .S(_13794_),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _16931_ (.A0(_13781_),
    .A1(\cpuregs[9][3] ),
    .S(_13794_),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_1 _16932_ (.A0(_13782_),
    .A1(\cpuregs[9][2] ),
    .S(_13794_),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_1 _16933_ (.A0(_13783_),
    .A1(\cpuregs[9][1] ),
    .S(_13789_),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_1 _16934_ (.A0(_13784_),
    .A1(\cpuregs[9][0] ),
    .S(_13789_),
    .X(_03664_));
 sky130_fd_sc_hd__o21ai_4 _16935_ (.A1(_12849_),
    .A2(_12842_),
    .B1(_12674_),
    .Y(_13795_));
 sky130_fd_sc_hd__buf_4 _16936_ (.A(_13795_),
    .X(_13796_));
 sky130_fd_sc_hd__mux2_1 _16937_ (.A0(_02467_),
    .A1(_12808_),
    .S(_13796_),
    .X(_03663_));
 sky130_fd_sc_hd__buf_4 _16938_ (.A(net361),
    .X(_13797_));
 sky130_fd_sc_hd__mux2_1 _16939_ (.A0(_02466_),
    .A1(_13797_),
    .S(_13796_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_4 _16940_ (.A(net359),
    .X(_13798_));
 sky130_fd_sc_hd__mux2_1 _16941_ (.A0(_02464_),
    .A1(_13798_),
    .S(_13796_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_4 _16942_ (.A(net358),
    .X(_13799_));
 sky130_fd_sc_hd__mux2_1 _16943_ (.A0(_02463_),
    .A1(_13799_),
    .S(_13796_),
    .X(_03660_));
 sky130_fd_sc_hd__clkbuf_4 _16944_ (.A(net357),
    .X(_13800_));
 sky130_fd_sc_hd__mux2_1 _16945_ (.A0(_02462_),
    .A1(_13800_),
    .S(_13796_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_4 _16946_ (.A(net356),
    .X(_13801_));
 sky130_fd_sc_hd__clkbuf_2 _16947_ (.A(_13795_),
    .X(_13802_));
 sky130_fd_sc_hd__buf_2 _16948_ (.A(_13802_),
    .X(_13803_));
 sky130_fd_sc_hd__mux2_1 _16949_ (.A0(_02461_),
    .A1(_13801_),
    .S(_13803_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_4 _16950_ (.A(net355),
    .X(_13804_));
 sky130_fd_sc_hd__mux2_1 _16951_ (.A0(_02460_),
    .A1(_13804_),
    .S(_13803_),
    .X(_03657_));
 sky130_fd_sc_hd__buf_6 _16952_ (.A(net354),
    .X(_13805_));
 sky130_fd_sc_hd__mux2_1 _16953_ (.A0(_02459_),
    .A1(_13805_),
    .S(_13803_),
    .X(_03656_));
 sky130_fd_sc_hd__buf_4 _16954_ (.A(net353),
    .X(_13806_));
 sky130_fd_sc_hd__mux2_1 _16955_ (.A0(_02458_),
    .A1(_13806_),
    .S(_13803_),
    .X(_03655_));
 sky130_fd_sc_hd__buf_4 _16956_ (.A(net352),
    .X(_13807_));
 sky130_fd_sc_hd__mux2_1 _16957_ (.A0(_02457_),
    .A1(_13807_),
    .S(_13803_),
    .X(_03654_));
 sky130_fd_sc_hd__buf_4 _16958_ (.A(net351),
    .X(_13808_));
 sky130_fd_sc_hd__mux2_1 _16959_ (.A0(_02456_),
    .A1(_13808_),
    .S(_13803_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_4 _16960_ (.A(net350),
    .X(_13809_));
 sky130_fd_sc_hd__buf_2 _16961_ (.A(_13802_),
    .X(_13810_));
 sky130_fd_sc_hd__mux2_1 _16962_ (.A0(_02455_),
    .A1(_13809_),
    .S(_13810_),
    .X(_03652_));
 sky130_fd_sc_hd__buf_4 _16963_ (.A(net348),
    .X(_13811_));
 sky130_fd_sc_hd__mux2_1 _16964_ (.A0(_02453_),
    .A1(_13811_),
    .S(_13810_),
    .X(_03651_));
 sky130_fd_sc_hd__buf_4 _16965_ (.A(net347),
    .X(_13812_));
 sky130_fd_sc_hd__mux2_1 _16966_ (.A0(_02452_),
    .A1(_13812_),
    .S(_13810_),
    .X(_03650_));
 sky130_fd_sc_hd__buf_4 _16967_ (.A(net346),
    .X(_13813_));
 sky130_fd_sc_hd__mux2_1 _16968_ (.A0(_02451_),
    .A1(_13813_),
    .S(_13810_),
    .X(_03649_));
 sky130_fd_sc_hd__buf_4 _16969_ (.A(net345),
    .X(_13814_));
 sky130_fd_sc_hd__mux2_1 _16970_ (.A0(_02450_),
    .A1(_13814_),
    .S(_13810_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_4 _16971_ (.A(net344),
    .X(_13815_));
 sky130_fd_sc_hd__mux2_1 _16972_ (.A0(_02449_),
    .A1(_13815_),
    .S(_13810_),
    .X(_03647_));
 sky130_fd_sc_hd__buf_4 _16973_ (.A(net343),
    .X(_13816_));
 sky130_fd_sc_hd__buf_2 _16974_ (.A(_13802_),
    .X(_13817_));
 sky130_fd_sc_hd__mux2_1 _16975_ (.A0(_02448_),
    .A1(_13816_),
    .S(_13817_),
    .X(_03646_));
 sky130_fd_sc_hd__buf_4 _16976_ (.A(net342),
    .X(_13818_));
 sky130_fd_sc_hd__mux2_1 _16977_ (.A0(_02447_),
    .A1(_13818_),
    .S(_13817_),
    .X(_03645_));
 sky130_fd_sc_hd__buf_4 _16978_ (.A(net341),
    .X(_13819_));
 sky130_fd_sc_hd__mux2_1 _16979_ (.A0(_02446_),
    .A1(_13819_),
    .S(_13817_),
    .X(_03644_));
 sky130_fd_sc_hd__buf_4 _16980_ (.A(net340),
    .X(_13820_));
 sky130_fd_sc_hd__mux2_1 _16981_ (.A0(_02445_),
    .A1(_13820_),
    .S(_13817_),
    .X(_03643_));
 sky130_fd_sc_hd__buf_4 _16982_ (.A(net339),
    .X(_13821_));
 sky130_fd_sc_hd__mux2_1 _16983_ (.A0(_02444_),
    .A1(_13821_),
    .S(_13817_),
    .X(_03642_));
 sky130_fd_sc_hd__buf_4 _16984_ (.A(net369),
    .X(_13822_));
 sky130_fd_sc_hd__mux2_1 _16985_ (.A0(_02474_),
    .A1(_13822_),
    .S(_13817_),
    .X(_03641_));
 sky130_fd_sc_hd__buf_4 _16986_ (.A(net368),
    .X(_13823_));
 sky130_fd_sc_hd__buf_2 _16987_ (.A(_13795_),
    .X(_13824_));
 sky130_fd_sc_hd__mux2_1 _16988_ (.A0(_02473_),
    .A1(_13823_),
    .S(_13824_),
    .X(_03640_));
 sky130_fd_sc_hd__buf_2 _16989_ (.A(net229),
    .X(_13825_));
 sky130_fd_sc_hd__buf_6 _16990_ (.A(_13825_),
    .X(_13826_));
 sky130_fd_sc_hd__mux2_1 _16991_ (.A0(_02472_),
    .A1(_13826_),
    .S(_13824_),
    .X(_03639_));
 sky130_fd_sc_hd__buf_2 _16992_ (.A(net228),
    .X(_13827_));
 sky130_fd_sc_hd__buf_6 _16993_ (.A(_13827_),
    .X(_13828_));
 sky130_fd_sc_hd__mux2_1 _16994_ (.A0(_02471_),
    .A1(_13828_),
    .S(_13824_),
    .X(_03638_));
 sky130_fd_sc_hd__clkbuf_4 _16995_ (.A(net227),
    .X(_13829_));
 sky130_fd_sc_hd__buf_4 _16996_ (.A(_13829_),
    .X(_13830_));
 sky130_fd_sc_hd__mux2_1 _16997_ (.A0(_02470_),
    .A1(_13830_),
    .S(_13824_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_2 _16998_ (.A(net226),
    .X(_13831_));
 sky130_fd_sc_hd__buf_4 _16999_ (.A(_13831_),
    .X(_13832_));
 sky130_fd_sc_hd__mux2_1 _17000_ (.A0(_02469_),
    .A1(_13832_),
    .S(_13824_),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_2 _17001_ (.A(net225),
    .X(_13833_));
 sky130_fd_sc_hd__buf_4 _17002_ (.A(_13833_),
    .X(_13834_));
 sky130_fd_sc_hd__mux2_1 _17003_ (.A0(_02468_),
    .A1(_13834_),
    .S(_13824_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_4 _17004_ (.A(net222),
    .X(_13835_));
 sky130_fd_sc_hd__buf_4 _17005_ (.A(_13835_),
    .X(_13836_));
 sky130_fd_sc_hd__mux2_1 _17006_ (.A0(_02465_),
    .A1(_13836_),
    .S(_13802_),
    .X(_03634_));
 sky130_fd_sc_hd__clkbuf_4 _17007_ (.A(net492),
    .X(_13837_));
 sky130_fd_sc_hd__buf_4 _17008_ (.A(_13837_),
    .X(_13838_));
 sky130_fd_sc_hd__mux2_1 _17009_ (.A0(_02454_),
    .A1(_13838_),
    .S(_13802_),
    .X(_03633_));
 sky130_fd_sc_hd__buf_4 _17010_ (.A(net200),
    .X(_13839_));
 sky130_fd_sc_hd__clkbuf_4 _17011_ (.A(_13839_),
    .X(_13840_));
 sky130_fd_sc_hd__mux2_1 _17012_ (.A0(_02443_),
    .A1(_13840_),
    .S(_13802_),
    .X(_03632_));
 sky130_fd_sc_hd__nand3b_4 _17013_ (.A_N(_13742_),
    .B(_13746_),
    .C(_13739_),
    .Y(_13841_));
 sky130_fd_sc_hd__buf_8 _17014_ (.A(_13841_),
    .X(_13842_));
 sky130_fd_sc_hd__buf_4 _17015_ (.A(_13842_),
    .X(_13843_));
 sky130_fd_sc_hd__mux2_1 _17016_ (.A0(_13734_),
    .A1(\cpuregs[4][31] ),
    .S(_13843_),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_1 _17017_ (.A0(_13750_),
    .A1(\cpuregs[4][30] ),
    .S(_13843_),
    .X(_03630_));
 sky130_fd_sc_hd__mux2_1 _17018_ (.A0(_13751_),
    .A1(\cpuregs[4][29] ),
    .S(_13843_),
    .X(_03629_));
 sky130_fd_sc_hd__mux2_1 _17019_ (.A0(_13752_),
    .A1(\cpuregs[4][28] ),
    .S(_13843_),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_1 _17020_ (.A0(_13753_),
    .A1(\cpuregs[4][27] ),
    .S(_13843_),
    .X(_03627_));
 sky130_fd_sc_hd__mux2_1 _17021_ (.A0(_13754_),
    .A1(\cpuregs[4][26] ),
    .S(_13843_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_4 _17022_ (.A(_13842_),
    .X(_13844_));
 sky130_fd_sc_hd__mux2_1 _17023_ (.A0(_13755_),
    .A1(\cpuregs[4][25] ),
    .S(_13844_),
    .X(_03625_));
 sky130_fd_sc_hd__mux2_1 _17024_ (.A0(_13757_),
    .A1(\cpuregs[4][24] ),
    .S(_13844_),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_1 _17025_ (.A0(_13758_),
    .A1(\cpuregs[4][23] ),
    .S(_13844_),
    .X(_03623_));
 sky130_fd_sc_hd__mux2_1 _17026_ (.A0(_13759_),
    .A1(\cpuregs[4][22] ),
    .S(_13844_),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_1 _17027_ (.A0(_13760_),
    .A1(\cpuregs[4][21] ),
    .S(_13844_),
    .X(_03621_));
 sky130_fd_sc_hd__mux2_1 _17028_ (.A0(_13761_),
    .A1(\cpuregs[4][20] ),
    .S(_13844_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_2 _17029_ (.A(_13842_),
    .X(_13845_));
 sky130_fd_sc_hd__mux2_1 _17030_ (.A0(_13762_),
    .A1(\cpuregs[4][19] ),
    .S(_13845_),
    .X(_03619_));
 sky130_fd_sc_hd__mux2_1 _17031_ (.A0(_13764_),
    .A1(\cpuregs[4][18] ),
    .S(_13845_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_1 _17032_ (.A0(_13765_),
    .A1(\cpuregs[4][17] ),
    .S(_13845_),
    .X(_03617_));
 sky130_fd_sc_hd__mux2_1 _17033_ (.A0(_13766_),
    .A1(\cpuregs[4][16] ),
    .S(_13845_),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _17034_ (.A0(_13767_),
    .A1(\cpuregs[4][15] ),
    .S(_13845_),
    .X(_03615_));
 sky130_fd_sc_hd__mux2_1 _17035_ (.A0(_13768_),
    .A1(\cpuregs[4][14] ),
    .S(_13845_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_4 _17036_ (.A(_13842_),
    .X(_13846_));
 sky130_fd_sc_hd__mux2_1 _17037_ (.A0(_13769_),
    .A1(\cpuregs[4][13] ),
    .S(_13846_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _17038_ (.A0(_13771_),
    .A1(\cpuregs[4][12] ),
    .S(_13846_),
    .X(_03612_));
 sky130_fd_sc_hd__mux2_1 _17039_ (.A0(_13772_),
    .A1(\cpuregs[4][11] ),
    .S(_13846_),
    .X(_03611_));
 sky130_fd_sc_hd__mux2_1 _17040_ (.A0(_13773_),
    .A1(\cpuregs[4][10] ),
    .S(_13846_),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _17041_ (.A0(_13774_),
    .A1(\cpuregs[4][9] ),
    .S(_13846_),
    .X(_03609_));
 sky130_fd_sc_hd__mux2_1 _17042_ (.A0(_13775_),
    .A1(\cpuregs[4][8] ),
    .S(_13846_),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_4 _17043_ (.A(_13841_),
    .X(_13847_));
 sky130_fd_sc_hd__mux2_1 _17044_ (.A0(_13776_),
    .A1(\cpuregs[4][7] ),
    .S(_13847_),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _17045_ (.A0(_13778_),
    .A1(\cpuregs[4][6] ),
    .S(_13847_),
    .X(_03606_));
 sky130_fd_sc_hd__mux2_1 _17046_ (.A0(_13779_),
    .A1(\cpuregs[4][5] ),
    .S(_13847_),
    .X(_03605_));
 sky130_fd_sc_hd__mux2_1 _17047_ (.A0(_13780_),
    .A1(\cpuregs[4][4] ),
    .S(_13847_),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_1 _17048_ (.A0(_13781_),
    .A1(\cpuregs[4][3] ),
    .S(_13847_),
    .X(_03603_));
 sky130_fd_sc_hd__mux2_1 _17049_ (.A0(_13782_),
    .A1(\cpuregs[4][2] ),
    .S(_13847_),
    .X(_03602_));
 sky130_fd_sc_hd__mux2_1 _17050_ (.A0(_13783_),
    .A1(\cpuregs[4][1] ),
    .S(_13842_),
    .X(_03601_));
 sky130_fd_sc_hd__mux2_1 _17051_ (.A0(_13784_),
    .A1(\cpuregs[4][0] ),
    .S(_13842_),
    .X(_03600_));
 sky130_fd_sc_hd__nor3b_4 _17052_ (.A(_13785_),
    .B(_13742_),
    .C_N(\latched_rd[1] ),
    .Y(_13848_));
 sky130_fd_sc_hd__nor3b_4 _17053_ (.A(_13745_),
    .B(_13744_),
    .C_N(\latched_rd[4] ),
    .Y(_13849_));
 sky130_fd_sc_hd__nand2_1 _17054_ (.A(_13848_),
    .B(_13849_),
    .Y(_13850_));
 sky130_fd_sc_hd__buf_6 _17055_ (.A(_13850_),
    .X(_13851_));
 sky130_fd_sc_hd__clkbuf_4 _17056_ (.A(_13851_),
    .X(_13852_));
 sky130_fd_sc_hd__mux2_1 _17057_ (.A0(_13734_),
    .A1(\cpuregs[19][31] ),
    .S(_13852_),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_1 _17058_ (.A0(_13750_),
    .A1(\cpuregs[19][30] ),
    .S(_13852_),
    .X(_03598_));
 sky130_fd_sc_hd__mux2_1 _17059_ (.A0(_13751_),
    .A1(\cpuregs[19][29] ),
    .S(_13852_),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_1 _17060_ (.A0(_13752_),
    .A1(\cpuregs[19][28] ),
    .S(_13852_),
    .X(_03596_));
 sky130_fd_sc_hd__mux2_1 _17061_ (.A0(_13753_),
    .A1(\cpuregs[19][27] ),
    .S(_13852_),
    .X(_03595_));
 sky130_fd_sc_hd__mux2_1 _17062_ (.A0(_13754_),
    .A1(\cpuregs[19][26] ),
    .S(_13852_),
    .X(_03594_));
 sky130_fd_sc_hd__buf_2 _17063_ (.A(_13851_),
    .X(_13853_));
 sky130_fd_sc_hd__mux2_1 _17064_ (.A0(_13755_),
    .A1(\cpuregs[19][25] ),
    .S(_13853_),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_1 _17065_ (.A0(_13757_),
    .A1(\cpuregs[19][24] ),
    .S(_13853_),
    .X(_03592_));
 sky130_fd_sc_hd__mux2_1 _17066_ (.A0(_13758_),
    .A1(\cpuregs[19][23] ),
    .S(_13853_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_1 _17067_ (.A0(_13759_),
    .A1(\cpuregs[19][22] ),
    .S(_13853_),
    .X(_03590_));
 sky130_fd_sc_hd__mux2_1 _17068_ (.A0(_13760_),
    .A1(\cpuregs[19][21] ),
    .S(_13853_),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_1 _17069_ (.A0(_13761_),
    .A1(\cpuregs[19][20] ),
    .S(_13853_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_4 _17070_ (.A(_13851_),
    .X(_13854_));
 sky130_fd_sc_hd__mux2_1 _17071_ (.A0(_13762_),
    .A1(\cpuregs[19][19] ),
    .S(_13854_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _17072_ (.A0(_13764_),
    .A1(\cpuregs[19][18] ),
    .S(_13854_),
    .X(_03586_));
 sky130_fd_sc_hd__mux2_1 _17073_ (.A0(_13765_),
    .A1(\cpuregs[19][17] ),
    .S(_13854_),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_1 _17074_ (.A0(_13766_),
    .A1(\cpuregs[19][16] ),
    .S(_13854_),
    .X(_03584_));
 sky130_fd_sc_hd__mux2_1 _17075_ (.A0(_13767_),
    .A1(\cpuregs[19][15] ),
    .S(_13854_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _17076_ (.A0(_13768_),
    .A1(\cpuregs[19][14] ),
    .S(_13854_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_4 _17077_ (.A(_13851_),
    .X(_13855_));
 sky130_fd_sc_hd__mux2_1 _17078_ (.A0(_13769_),
    .A1(\cpuregs[19][13] ),
    .S(_13855_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_1 _17079_ (.A0(_13771_),
    .A1(\cpuregs[19][12] ),
    .S(_13855_),
    .X(_03580_));
 sky130_fd_sc_hd__mux2_1 _17080_ (.A0(_13772_),
    .A1(\cpuregs[19][11] ),
    .S(_13855_),
    .X(_03579_));
 sky130_fd_sc_hd__mux2_1 _17081_ (.A0(_13773_),
    .A1(\cpuregs[19][10] ),
    .S(_13855_),
    .X(_03578_));
 sky130_fd_sc_hd__mux2_1 _17082_ (.A0(_13774_),
    .A1(\cpuregs[19][9] ),
    .S(_13855_),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_1 _17083_ (.A0(_13775_),
    .A1(\cpuregs[19][8] ),
    .S(_13855_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_4 _17084_ (.A(_13850_),
    .X(_13856_));
 sky130_fd_sc_hd__mux2_1 _17085_ (.A0(_13776_),
    .A1(\cpuregs[19][7] ),
    .S(_13856_),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_1 _17086_ (.A0(_13778_),
    .A1(\cpuregs[19][6] ),
    .S(_13856_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_1 _17087_ (.A0(_13779_),
    .A1(\cpuregs[19][5] ),
    .S(_13856_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _17088_ (.A0(_13780_),
    .A1(\cpuregs[19][4] ),
    .S(_13856_),
    .X(_03572_));
 sky130_fd_sc_hd__mux2_1 _17089_ (.A0(_13781_),
    .A1(\cpuregs[19][3] ),
    .S(_13856_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_1 _17090_ (.A0(_13782_),
    .A1(\cpuregs[19][2] ),
    .S(_13856_),
    .X(_03570_));
 sky130_fd_sc_hd__mux2_1 _17091_ (.A0(_13783_),
    .A1(\cpuregs[19][1] ),
    .S(_13851_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _17092_ (.A0(_13784_),
    .A1(\cpuregs[19][0] ),
    .S(_13851_),
    .X(_03568_));
 sky130_fd_sc_hd__nand3_4 _17093_ (.A(_12665_),
    .B(_12678_),
    .C(_12638_),
    .Y(_13857_));
 sky130_fd_sc_hd__nand3b_4 _17094_ (.A_N(_13857_),
    .B(_12976_),
    .C(_12669_),
    .Y(_13858_));
 sky130_fd_sc_hd__clkbuf_4 _17095_ (.A(_13858_),
    .X(_13859_));
 sky130_fd_sc_hd__clkbuf_8 _17096_ (.A(_13859_),
    .X(_13860_));
 sky130_fd_sc_hd__mux2_1 _17097_ (.A0(net224),
    .A1(net262),
    .S(_13860_),
    .X(_03567_));
 sky130_fd_sc_hd__mux2_1 _17098_ (.A0(net223),
    .A1(net261),
    .S(_13860_),
    .X(_03566_));
 sky130_fd_sc_hd__mux2_1 _17099_ (.A0(net221),
    .A1(net259),
    .S(_13860_),
    .X(_03565_));
 sky130_fd_sc_hd__mux2_1 _17100_ (.A0(net220),
    .A1(net258),
    .S(_13860_),
    .X(_03564_));
 sky130_fd_sc_hd__mux2_1 _17101_ (.A0(net219),
    .A1(net257),
    .S(_13860_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _17102_ (.A0(net218),
    .A1(net256),
    .S(_13860_),
    .X(_03562_));
 sky130_fd_sc_hd__buf_6 _17103_ (.A(_13859_),
    .X(_13861_));
 sky130_fd_sc_hd__mux2_1 _17104_ (.A0(net217),
    .A1(net255),
    .S(_13861_),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _17105_ (.A0(net216),
    .A1(net254),
    .S(_13861_),
    .X(_03560_));
 sky130_fd_sc_hd__mux2_1 _17106_ (.A0(net215),
    .A1(net253),
    .S(_13861_),
    .X(_03559_));
 sky130_fd_sc_hd__mux2_1 _17107_ (.A0(net214),
    .A1(net252),
    .S(_13861_),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_1 _17108_ (.A0(net213),
    .A1(net251),
    .S(_13861_),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_1 _17109_ (.A0(net212),
    .A1(net250),
    .S(_13861_),
    .X(_03556_));
 sky130_fd_sc_hd__buf_8 _17110_ (.A(_13859_),
    .X(_13862_));
 sky130_fd_sc_hd__mux2_1 _17111_ (.A0(net210),
    .A1(net248),
    .S(_13862_),
    .X(_03555_));
 sky130_fd_sc_hd__mux2_1 _17112_ (.A0(net209),
    .A1(net247),
    .S(_13862_),
    .X(_03554_));
 sky130_fd_sc_hd__mux2_1 _17113_ (.A0(net208),
    .A1(net246),
    .S(net423),
    .X(_03553_));
 sky130_fd_sc_hd__mux2_1 _17114_ (.A0(net207),
    .A1(net245),
    .S(net423),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _17115_ (.A0(net206),
    .A1(net244),
    .S(_13862_),
    .X(_03551_));
 sky130_fd_sc_hd__mux2_1 _17116_ (.A0(net205),
    .A1(net243),
    .S(_13862_),
    .X(_03550_));
 sky130_fd_sc_hd__buf_6 _17117_ (.A(_13859_),
    .X(_13863_));
 sky130_fd_sc_hd__mux2_1 _17118_ (.A0(net204),
    .A1(net242),
    .S(net422),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_1 _17119_ (.A0(net203),
    .A1(net241),
    .S(_13863_),
    .X(_03548_));
 sky130_fd_sc_hd__mux2_1 _17120_ (.A0(net202),
    .A1(net240),
    .S(_13863_),
    .X(_03547_));
 sky130_fd_sc_hd__mux2_1 _17121_ (.A0(net201),
    .A1(net239),
    .S(_13863_),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_1 _17122_ (.A0(net231),
    .A1(net269),
    .S(net422),
    .X(_03545_));
 sky130_fd_sc_hd__mux2_1 _17123_ (.A0(net230),
    .A1(net268),
    .S(net422),
    .X(_03544_));
 sky130_fd_sc_hd__buf_4 _17124_ (.A(_13858_),
    .X(_13864_));
 sky130_fd_sc_hd__mux2_1 _17125_ (.A0(_13826_),
    .A1(net267),
    .S(_13864_),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_1 _17126_ (.A0(_13828_),
    .A1(net266),
    .S(_13864_),
    .X(_03542_));
 sky130_fd_sc_hd__mux2_1 _17127_ (.A0(_13830_),
    .A1(net265),
    .S(_13864_),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_1 _17128_ (.A0(_13832_),
    .A1(net264),
    .S(_13864_),
    .X(_03540_));
 sky130_fd_sc_hd__mux2_1 _17129_ (.A0(_13834_),
    .A1(net263),
    .S(_13864_),
    .X(_03539_));
 sky130_fd_sc_hd__mux2_1 _17130_ (.A0(_13836_),
    .A1(net260),
    .S(_13864_),
    .X(_03538_));
 sky130_fd_sc_hd__mux2_1 _17131_ (.A0(_13838_),
    .A1(net249),
    .S(_13859_),
    .X(_03537_));
 sky130_fd_sc_hd__mux2_1 _17132_ (.A0(_13840_),
    .A1(net238),
    .S(_13859_),
    .X(_03536_));
 sky130_fd_sc_hd__nand2_2 _17133_ (.A(_13848_),
    .B(_13746_),
    .Y(_13865_));
 sky130_fd_sc_hd__buf_8 _17134_ (.A(_13865_),
    .X(_13866_));
 sky130_fd_sc_hd__buf_4 _17135_ (.A(_13866_),
    .X(_13867_));
 sky130_fd_sc_hd__mux2_1 _17136_ (.A0(_13734_),
    .A1(\cpuregs[7][31] ),
    .S(_13867_),
    .X(_03535_));
 sky130_fd_sc_hd__mux2_1 _17137_ (.A0(_13750_),
    .A1(\cpuregs[7][30] ),
    .S(_13867_),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_1 _17138_ (.A0(_13751_),
    .A1(\cpuregs[7][29] ),
    .S(_13867_),
    .X(_03533_));
 sky130_fd_sc_hd__mux2_1 _17139_ (.A0(_13752_),
    .A1(\cpuregs[7][28] ),
    .S(_13867_),
    .X(_03532_));
 sky130_fd_sc_hd__mux2_1 _17140_ (.A0(_13753_),
    .A1(\cpuregs[7][27] ),
    .S(_13867_),
    .X(_03531_));
 sky130_fd_sc_hd__mux2_1 _17141_ (.A0(_13754_),
    .A1(\cpuregs[7][26] ),
    .S(_13867_),
    .X(_03530_));
 sky130_fd_sc_hd__buf_2 _17142_ (.A(_13866_),
    .X(_13868_));
 sky130_fd_sc_hd__mux2_1 _17143_ (.A0(_13755_),
    .A1(\cpuregs[7][25] ),
    .S(_13868_),
    .X(_03529_));
 sky130_fd_sc_hd__mux2_1 _17144_ (.A0(_13757_),
    .A1(\cpuregs[7][24] ),
    .S(_13868_),
    .X(_03528_));
 sky130_fd_sc_hd__mux2_1 _17145_ (.A0(_13758_),
    .A1(\cpuregs[7][23] ),
    .S(_13868_),
    .X(_03527_));
 sky130_fd_sc_hd__mux2_1 _17146_ (.A0(_13759_),
    .A1(\cpuregs[7][22] ),
    .S(_13868_),
    .X(_03526_));
 sky130_fd_sc_hd__mux2_1 _17147_ (.A0(_13760_),
    .A1(\cpuregs[7][21] ),
    .S(_13868_),
    .X(_03525_));
 sky130_fd_sc_hd__mux2_1 _17148_ (.A0(_13761_),
    .A1(\cpuregs[7][20] ),
    .S(_13868_),
    .X(_03524_));
 sky130_fd_sc_hd__buf_2 _17149_ (.A(_13866_),
    .X(_13869_));
 sky130_fd_sc_hd__mux2_1 _17150_ (.A0(_13762_),
    .A1(\cpuregs[7][19] ),
    .S(_13869_),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_1 _17151_ (.A0(_13764_),
    .A1(\cpuregs[7][18] ),
    .S(_13869_),
    .X(_03522_));
 sky130_fd_sc_hd__mux2_1 _17152_ (.A0(_13765_),
    .A1(\cpuregs[7][17] ),
    .S(_13869_),
    .X(_03521_));
 sky130_fd_sc_hd__mux2_1 _17153_ (.A0(_13766_),
    .A1(\cpuregs[7][16] ),
    .S(_13869_),
    .X(_03520_));
 sky130_fd_sc_hd__mux2_1 _17154_ (.A0(_13767_),
    .A1(\cpuregs[7][15] ),
    .S(_13869_),
    .X(_03519_));
 sky130_fd_sc_hd__mux2_1 _17155_ (.A0(_13768_),
    .A1(\cpuregs[7][14] ),
    .S(_13869_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_4 _17156_ (.A(_13866_),
    .X(_13870_));
 sky130_fd_sc_hd__mux2_1 _17157_ (.A0(_13769_),
    .A1(\cpuregs[7][13] ),
    .S(_13870_),
    .X(_03517_));
 sky130_fd_sc_hd__mux2_1 _17158_ (.A0(_13771_),
    .A1(\cpuregs[7][12] ),
    .S(_13870_),
    .X(_03516_));
 sky130_fd_sc_hd__mux2_1 _17159_ (.A0(_13772_),
    .A1(\cpuregs[7][11] ),
    .S(_13870_),
    .X(_03515_));
 sky130_fd_sc_hd__mux2_1 _17160_ (.A0(_13773_),
    .A1(\cpuregs[7][10] ),
    .S(_13870_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_1 _17161_ (.A0(_13774_),
    .A1(\cpuregs[7][9] ),
    .S(_13870_),
    .X(_03513_));
 sky130_fd_sc_hd__mux2_1 _17162_ (.A0(_13775_),
    .A1(\cpuregs[7][8] ),
    .S(_13870_),
    .X(_03512_));
 sky130_fd_sc_hd__clkbuf_4 _17163_ (.A(_13865_),
    .X(_13871_));
 sky130_fd_sc_hd__mux2_1 _17164_ (.A0(_13776_),
    .A1(\cpuregs[7][7] ),
    .S(_13871_),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_1 _17165_ (.A0(_13778_),
    .A1(\cpuregs[7][6] ),
    .S(_13871_),
    .X(_03510_));
 sky130_fd_sc_hd__mux2_1 _17166_ (.A0(_13779_),
    .A1(\cpuregs[7][5] ),
    .S(_13871_),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_1 _17167_ (.A0(_13780_),
    .A1(\cpuregs[7][4] ),
    .S(_13871_),
    .X(_03508_));
 sky130_fd_sc_hd__mux2_1 _17168_ (.A0(_13781_),
    .A1(\cpuregs[7][3] ),
    .S(_13871_),
    .X(_03507_));
 sky130_fd_sc_hd__mux2_1 _17169_ (.A0(_13782_),
    .A1(\cpuregs[7][2] ),
    .S(_13871_),
    .X(_03506_));
 sky130_fd_sc_hd__mux2_1 _17170_ (.A0(_13783_),
    .A1(\cpuregs[7][1] ),
    .S(_13866_),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_1 _17171_ (.A0(_13784_),
    .A1(\cpuregs[7][0] ),
    .S(_13866_),
    .X(_03504_));
 sky130_fd_sc_hd__buf_2 _17172_ (.A(_12852_),
    .X(_13872_));
 sky130_fd_sc_hd__and2b_1 _17173_ (.A_N(_00331_),
    .B(_12674_),
    .X(_13873_));
 sky130_fd_sc_hd__nor3b_1 _17174_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(_12846_),
    .C_N(\cpu_state[4] ),
    .Y(_13874_));
 sky130_vsdinv _17175_ (.A(_13874_),
    .Y(_13875_));
 sky130_fd_sc_hd__o211ai_2 _17176_ (.A1(instr_setq),
    .A2(_13872_),
    .B1(_13873_),
    .C1(_13875_),
    .Y(_13876_));
 sky130_fd_sc_hd__mux2_1 _17177_ (.A0(_15206_),
    .A1(\latched_rd[4] ),
    .S(_13876_),
    .X(_03503_));
 sky130_fd_sc_hd__nand3b_1 _17178_ (.A_N(\latched_rd[4] ),
    .B(_13745_),
    .C(_13744_),
    .Y(_13877_));
 sky130_vsdinv _17179_ (.A(_13877_),
    .Y(_13878_));
 sky130_fd_sc_hd__nand2_1 _17180_ (.A(_13848_),
    .B(_13878_),
    .Y(_13879_));
 sky130_fd_sc_hd__buf_6 _17181_ (.A(_13879_),
    .X(_13880_));
 sky130_fd_sc_hd__clkbuf_4 _17182_ (.A(_13880_),
    .X(_13881_));
 sky130_fd_sc_hd__mux2_1 _17183_ (.A0(_13734_),
    .A1(\cpuregs[15][31] ),
    .S(_13881_),
    .X(_03502_));
 sky130_fd_sc_hd__mux2_1 _17184_ (.A0(_13750_),
    .A1(\cpuregs[15][30] ),
    .S(_13881_),
    .X(_03501_));
 sky130_fd_sc_hd__mux2_1 _17185_ (.A0(_13751_),
    .A1(\cpuregs[15][29] ),
    .S(_13881_),
    .X(_03500_));
 sky130_fd_sc_hd__mux2_1 _17186_ (.A0(_13752_),
    .A1(\cpuregs[15][28] ),
    .S(_13881_),
    .X(_03499_));
 sky130_fd_sc_hd__mux2_1 _17187_ (.A0(_13753_),
    .A1(\cpuregs[15][27] ),
    .S(_13881_),
    .X(_03498_));
 sky130_fd_sc_hd__mux2_1 _17188_ (.A0(_13754_),
    .A1(\cpuregs[15][26] ),
    .S(_13881_),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_4 _17189_ (.A(_13880_),
    .X(_13882_));
 sky130_fd_sc_hd__mux2_1 _17190_ (.A0(_13755_),
    .A1(\cpuregs[15][25] ),
    .S(_13882_),
    .X(_03496_));
 sky130_fd_sc_hd__mux2_1 _17191_ (.A0(_13757_),
    .A1(\cpuregs[15][24] ),
    .S(_13882_),
    .X(_03495_));
 sky130_fd_sc_hd__mux2_1 _17192_ (.A0(_13758_),
    .A1(\cpuregs[15][23] ),
    .S(_13882_),
    .X(_03494_));
 sky130_fd_sc_hd__mux2_1 _17193_ (.A0(_13759_),
    .A1(\cpuregs[15][22] ),
    .S(_13882_),
    .X(_03493_));
 sky130_fd_sc_hd__mux2_1 _17194_ (.A0(_13760_),
    .A1(\cpuregs[15][21] ),
    .S(_13882_),
    .X(_03492_));
 sky130_fd_sc_hd__mux2_1 _17195_ (.A0(_13761_),
    .A1(\cpuregs[15][20] ),
    .S(_13882_),
    .X(_03491_));
 sky130_fd_sc_hd__clkbuf_4 _17196_ (.A(_13880_),
    .X(_13883_));
 sky130_fd_sc_hd__mux2_1 _17197_ (.A0(_13762_),
    .A1(\cpuregs[15][19] ),
    .S(_13883_),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_1 _17198_ (.A0(_13764_),
    .A1(\cpuregs[15][18] ),
    .S(_13883_),
    .X(_03489_));
 sky130_fd_sc_hd__mux2_1 _17199_ (.A0(_13765_),
    .A1(\cpuregs[15][17] ),
    .S(_13883_),
    .X(_03488_));
 sky130_fd_sc_hd__mux2_1 _17200_ (.A0(_13766_),
    .A1(\cpuregs[15][16] ),
    .S(_13883_),
    .X(_03487_));
 sky130_fd_sc_hd__mux2_1 _17201_ (.A0(_13767_),
    .A1(\cpuregs[15][15] ),
    .S(_13883_),
    .X(_03486_));
 sky130_fd_sc_hd__mux2_1 _17202_ (.A0(_13768_),
    .A1(\cpuregs[15][14] ),
    .S(_13883_),
    .X(_03485_));
 sky130_fd_sc_hd__clkbuf_4 _17203_ (.A(_13880_),
    .X(_13884_));
 sky130_fd_sc_hd__mux2_1 _17204_ (.A0(_13769_),
    .A1(\cpuregs[15][13] ),
    .S(_13884_),
    .X(_03484_));
 sky130_fd_sc_hd__mux2_1 _17205_ (.A0(_13771_),
    .A1(\cpuregs[15][12] ),
    .S(_13884_),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_1 _17206_ (.A0(_13772_),
    .A1(\cpuregs[15][11] ),
    .S(_13884_),
    .X(_03482_));
 sky130_fd_sc_hd__mux2_1 _17207_ (.A0(_13773_),
    .A1(\cpuregs[15][10] ),
    .S(_13884_),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_1 _17208_ (.A0(_13774_),
    .A1(\cpuregs[15][9] ),
    .S(_13884_),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_1 _17209_ (.A0(_13775_),
    .A1(\cpuregs[15][8] ),
    .S(_13884_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_4 _17210_ (.A(_13879_),
    .X(_13885_));
 sky130_fd_sc_hd__mux2_1 _17211_ (.A0(_13776_),
    .A1(\cpuregs[15][7] ),
    .S(_13885_),
    .X(_03478_));
 sky130_fd_sc_hd__mux2_1 _17212_ (.A0(_13778_),
    .A1(\cpuregs[15][6] ),
    .S(_13885_),
    .X(_03477_));
 sky130_fd_sc_hd__mux2_1 _17213_ (.A0(_13779_),
    .A1(\cpuregs[15][5] ),
    .S(_13885_),
    .X(_03476_));
 sky130_fd_sc_hd__mux2_1 _17214_ (.A0(_13780_),
    .A1(\cpuregs[15][4] ),
    .S(_13885_),
    .X(_03475_));
 sky130_fd_sc_hd__mux2_1 _17215_ (.A0(_13781_),
    .A1(\cpuregs[15][3] ),
    .S(_13885_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_1 _17216_ (.A0(_13782_),
    .A1(\cpuregs[15][2] ),
    .S(_13885_),
    .X(_03473_));
 sky130_fd_sc_hd__mux2_1 _17217_ (.A0(_13783_),
    .A1(\cpuregs[15][1] ),
    .S(_13880_),
    .X(_03472_));
 sky130_fd_sc_hd__mux2_1 _17218_ (.A0(_13784_),
    .A1(\cpuregs[15][0] ),
    .S(_13880_),
    .X(_03471_));
 sky130_fd_sc_hd__buf_1 _17219_ (.A(\cpuregs_wrdata[31] ),
    .X(_13886_));
 sky130_fd_sc_hd__nand2_1 _17220_ (.A(_13848_),
    .B(_13787_),
    .Y(_13887_));
 sky130_fd_sc_hd__buf_6 _17221_ (.A(_13887_),
    .X(_13888_));
 sky130_fd_sc_hd__clkbuf_4 _17222_ (.A(_13888_),
    .X(_13889_));
 sky130_fd_sc_hd__mux2_1 _17223_ (.A0(_13886_),
    .A1(\cpuregs[11][31] ),
    .S(_13889_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_2 _17224_ (.A(\cpuregs_wrdata[30] ),
    .X(_13890_));
 sky130_fd_sc_hd__mux2_1 _17225_ (.A0(_13890_),
    .A1(\cpuregs[11][30] ),
    .S(_13889_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_2 _17226_ (.A(\cpuregs_wrdata[29] ),
    .X(_13891_));
 sky130_fd_sc_hd__mux2_1 _17227_ (.A0(_13891_),
    .A1(\cpuregs[11][29] ),
    .S(_13889_),
    .X(_03468_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17228_ (.A(\cpuregs_wrdata[28] ),
    .X(_13892_));
 sky130_fd_sc_hd__mux2_1 _17229_ (.A0(_13892_),
    .A1(\cpuregs[11][28] ),
    .S(_13889_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_2 _17230_ (.A(\cpuregs_wrdata[27] ),
    .X(_13893_));
 sky130_fd_sc_hd__mux2_1 _17231_ (.A0(_13893_),
    .A1(\cpuregs[11][27] ),
    .S(_13889_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_2 _17232_ (.A(\cpuregs_wrdata[26] ),
    .X(_13894_));
 sky130_fd_sc_hd__mux2_1 _17233_ (.A0(_13894_),
    .A1(\cpuregs[11][26] ),
    .S(_13889_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_2 _17234_ (.A(\cpuregs_wrdata[25] ),
    .X(_13895_));
 sky130_fd_sc_hd__clkbuf_4 _17235_ (.A(_13888_),
    .X(_13896_));
 sky130_fd_sc_hd__mux2_1 _17236_ (.A0(_13895_),
    .A1(\cpuregs[11][25] ),
    .S(_13896_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_2 _17237_ (.A(\cpuregs_wrdata[24] ),
    .X(_13897_));
 sky130_fd_sc_hd__mux2_1 _17238_ (.A0(_13897_),
    .A1(\cpuregs[11][24] ),
    .S(_13896_),
    .X(_03463_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17239_ (.A(\cpuregs_wrdata[23] ),
    .X(_13898_));
 sky130_fd_sc_hd__mux2_1 _17240_ (.A0(_13898_),
    .A1(\cpuregs[11][23] ),
    .S(_13896_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_2 _17241_ (.A(\cpuregs_wrdata[22] ),
    .X(_13899_));
 sky130_fd_sc_hd__mux2_1 _17242_ (.A0(_13899_),
    .A1(\cpuregs[11][22] ),
    .S(_13896_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_2 _17243_ (.A(\cpuregs_wrdata[21] ),
    .X(_13900_));
 sky130_fd_sc_hd__mux2_1 _17244_ (.A0(_13900_),
    .A1(\cpuregs[11][21] ),
    .S(_13896_),
    .X(_03460_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17245_ (.A(\cpuregs_wrdata[20] ),
    .X(_13901_));
 sky130_fd_sc_hd__mux2_1 _17246_ (.A0(_13901_),
    .A1(\cpuregs[11][20] ),
    .S(_13896_),
    .X(_03459_));
 sky130_fd_sc_hd__clkbuf_2 _17247_ (.A(\cpuregs_wrdata[19] ),
    .X(_13902_));
 sky130_fd_sc_hd__clkbuf_4 _17248_ (.A(_13888_),
    .X(_13903_));
 sky130_fd_sc_hd__mux2_1 _17249_ (.A0(_13902_),
    .A1(\cpuregs[11][19] ),
    .S(_13903_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_2 _17250_ (.A(\cpuregs_wrdata[18] ),
    .X(_13904_));
 sky130_fd_sc_hd__mux2_1 _17251_ (.A0(_13904_),
    .A1(\cpuregs[11][18] ),
    .S(_13903_),
    .X(_03457_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17252_ (.A(\cpuregs_wrdata[17] ),
    .X(_13905_));
 sky130_fd_sc_hd__mux2_1 _17253_ (.A0(_13905_),
    .A1(\cpuregs[11][17] ),
    .S(_13903_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_2 _17254_ (.A(\cpuregs_wrdata[16] ),
    .X(_13906_));
 sky130_fd_sc_hd__mux2_1 _17255_ (.A0(_13906_),
    .A1(\cpuregs[11][16] ),
    .S(_13903_),
    .X(_03455_));
 sky130_fd_sc_hd__buf_1 _17256_ (.A(\cpuregs_wrdata[15] ),
    .X(_13907_));
 sky130_fd_sc_hd__mux2_1 _17257_ (.A0(_13907_),
    .A1(\cpuregs[11][15] ),
    .S(_13903_),
    .X(_03454_));
 sky130_fd_sc_hd__buf_1 _17258_ (.A(\cpuregs_wrdata[14] ),
    .X(_13908_));
 sky130_fd_sc_hd__mux2_1 _17259_ (.A0(_13908_),
    .A1(\cpuregs[11][14] ),
    .S(_13903_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_2 _17260_ (.A(\cpuregs_wrdata[13] ),
    .X(_13909_));
 sky130_fd_sc_hd__clkbuf_4 _17261_ (.A(_13888_),
    .X(_13910_));
 sky130_fd_sc_hd__mux2_1 _17262_ (.A0(_13909_),
    .A1(\cpuregs[11][13] ),
    .S(_13910_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_2 _17263_ (.A(\cpuregs_wrdata[12] ),
    .X(_13911_));
 sky130_fd_sc_hd__mux2_1 _17264_ (.A0(_13911_),
    .A1(\cpuregs[11][12] ),
    .S(_13910_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_2 _17265_ (.A(\cpuregs_wrdata[11] ),
    .X(_13912_));
 sky130_fd_sc_hd__mux2_1 _17266_ (.A0(_13912_),
    .A1(\cpuregs[11][11] ),
    .S(_13910_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_2 _17267_ (.A(\cpuregs_wrdata[10] ),
    .X(_13913_));
 sky130_fd_sc_hd__mux2_1 _17268_ (.A0(_13913_),
    .A1(\cpuregs[11][10] ),
    .S(_13910_),
    .X(_03449_));
 sky130_fd_sc_hd__buf_1 _17269_ (.A(\cpuregs_wrdata[9] ),
    .X(_13914_));
 sky130_fd_sc_hd__mux2_1 _17270_ (.A0(_13914_),
    .A1(\cpuregs[11][9] ),
    .S(_13910_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_2 _17271_ (.A(\cpuregs_wrdata[8] ),
    .X(_13915_));
 sky130_fd_sc_hd__mux2_1 _17272_ (.A0(_13915_),
    .A1(\cpuregs[11][8] ),
    .S(_13910_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_2 _17273_ (.A(\cpuregs_wrdata[7] ),
    .X(_13916_));
 sky130_fd_sc_hd__clkbuf_4 _17274_ (.A(_13887_),
    .X(_13917_));
 sky130_fd_sc_hd__mux2_1 _17275_ (.A0(_13916_),
    .A1(\cpuregs[11][7] ),
    .S(_13917_),
    .X(_03446_));
 sky130_fd_sc_hd__clkbuf_2 _17276_ (.A(\cpuregs_wrdata[6] ),
    .X(_13918_));
 sky130_fd_sc_hd__mux2_1 _17277_ (.A0(_13918_),
    .A1(\cpuregs[11][6] ),
    .S(_13917_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_2 _17278_ (.A(\cpuregs_wrdata[5] ),
    .X(_13919_));
 sky130_fd_sc_hd__mux2_1 _17279_ (.A0(_13919_),
    .A1(\cpuregs[11][5] ),
    .S(_13917_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_2 _17280_ (.A(\cpuregs_wrdata[4] ),
    .X(_13920_));
 sky130_fd_sc_hd__mux2_1 _17281_ (.A0(_13920_),
    .A1(\cpuregs[11][4] ),
    .S(_13917_),
    .X(_03443_));
 sky130_fd_sc_hd__clkbuf_2 _17282_ (.A(\cpuregs_wrdata[3] ),
    .X(_13921_));
 sky130_fd_sc_hd__mux2_1 _17283_ (.A0(_13921_),
    .A1(\cpuregs[11][3] ),
    .S(_13917_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_2 _17284_ (.A(\cpuregs_wrdata[2] ),
    .X(_13922_));
 sky130_fd_sc_hd__mux2_1 _17285_ (.A0(_13922_),
    .A1(\cpuregs[11][2] ),
    .S(_13917_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_2 _17286_ (.A(\cpuregs_wrdata[1] ),
    .X(_13923_));
 sky130_fd_sc_hd__mux2_1 _17287_ (.A0(_13923_),
    .A1(\cpuregs[11][1] ),
    .S(_13888_),
    .X(_03440_));
 sky130_fd_sc_hd__buf_1 _17288_ (.A(\cpuregs_wrdata[0] ),
    .X(_13924_));
 sky130_fd_sc_hd__mux2_1 _17289_ (.A0(_13924_),
    .A1(\cpuregs[11][0] ),
    .S(_13888_),
    .X(_03439_));
 sky130_fd_sc_hd__nand2_1 _17290_ (.A(_13848_),
    .B(_13738_),
    .Y(_13925_));
 sky130_fd_sc_hd__buf_6 _17291_ (.A(_13925_),
    .X(_13926_));
 sky130_fd_sc_hd__buf_4 _17292_ (.A(_13926_),
    .X(_13927_));
 sky130_fd_sc_hd__mux2_1 _17293_ (.A0(_13886_),
    .A1(\cpuregs[3][31] ),
    .S(_13927_),
    .X(_03438_));
 sky130_fd_sc_hd__mux2_1 _17294_ (.A0(_13890_),
    .A1(\cpuregs[3][30] ),
    .S(_13927_),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_1 _17295_ (.A0(_13891_),
    .A1(\cpuregs[3][29] ),
    .S(_13927_),
    .X(_03436_));
 sky130_fd_sc_hd__mux2_1 _17296_ (.A0(_13892_),
    .A1(\cpuregs[3][28] ),
    .S(_13927_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _17297_ (.A0(_13893_),
    .A1(\cpuregs[3][27] ),
    .S(_13927_),
    .X(_03434_));
 sky130_fd_sc_hd__mux2_1 _17298_ (.A0(_13894_),
    .A1(\cpuregs[3][26] ),
    .S(_13927_),
    .X(_03433_));
 sky130_fd_sc_hd__clkbuf_4 _17299_ (.A(_13926_),
    .X(_13928_));
 sky130_fd_sc_hd__mux2_1 _17300_ (.A0(_13895_),
    .A1(\cpuregs[3][25] ),
    .S(_13928_),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_1 _17301_ (.A0(_13897_),
    .A1(\cpuregs[3][24] ),
    .S(_13928_),
    .X(_03431_));
 sky130_fd_sc_hd__mux2_1 _17302_ (.A0(_13898_),
    .A1(\cpuregs[3][23] ),
    .S(_13928_),
    .X(_03430_));
 sky130_fd_sc_hd__mux2_1 _17303_ (.A0(_13899_),
    .A1(\cpuregs[3][22] ),
    .S(_13928_),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_1 _17304_ (.A0(_13900_),
    .A1(\cpuregs[3][21] ),
    .S(_13928_),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_1 _17305_ (.A0(_13901_),
    .A1(\cpuregs[3][20] ),
    .S(_13928_),
    .X(_03427_));
 sky130_fd_sc_hd__clkbuf_4 _17306_ (.A(_13926_),
    .X(_13929_));
 sky130_fd_sc_hd__mux2_1 _17307_ (.A0(_13902_),
    .A1(\cpuregs[3][19] ),
    .S(_13929_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _17308_ (.A0(_13904_),
    .A1(\cpuregs[3][18] ),
    .S(_13929_),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_1 _17309_ (.A0(_13905_),
    .A1(\cpuregs[3][17] ),
    .S(_13929_),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_1 _17310_ (.A0(_13906_),
    .A1(\cpuregs[3][16] ),
    .S(_13929_),
    .X(_03423_));
 sky130_fd_sc_hd__mux2_1 _17311_ (.A0(_13907_),
    .A1(\cpuregs[3][15] ),
    .S(_13929_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_1 _17312_ (.A0(_13908_),
    .A1(\cpuregs[3][14] ),
    .S(_13929_),
    .X(_03421_));
 sky130_fd_sc_hd__buf_4 _17313_ (.A(_13926_),
    .X(_13930_));
 sky130_fd_sc_hd__mux2_1 _17314_ (.A0(_13909_),
    .A1(\cpuregs[3][13] ),
    .S(_13930_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _17315_ (.A0(_13911_),
    .A1(\cpuregs[3][12] ),
    .S(_13930_),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_1 _17316_ (.A0(_13912_),
    .A1(\cpuregs[3][11] ),
    .S(_13930_),
    .X(_03418_));
 sky130_fd_sc_hd__mux2_1 _17317_ (.A0(_13913_),
    .A1(\cpuregs[3][10] ),
    .S(_13930_),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_1 _17318_ (.A0(_13914_),
    .A1(\cpuregs[3][9] ),
    .S(_13930_),
    .X(_03416_));
 sky130_fd_sc_hd__mux2_1 _17319_ (.A0(_13915_),
    .A1(\cpuregs[3][8] ),
    .S(_13930_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_4 _17320_ (.A(_13925_),
    .X(_13931_));
 sky130_fd_sc_hd__mux2_1 _17321_ (.A0(_13916_),
    .A1(\cpuregs[3][7] ),
    .S(_13931_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _17322_ (.A0(_13918_),
    .A1(\cpuregs[3][6] ),
    .S(_13931_),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_1 _17323_ (.A0(_13919_),
    .A1(\cpuregs[3][5] ),
    .S(_13931_),
    .X(_03412_));
 sky130_fd_sc_hd__mux2_1 _17324_ (.A0(_13920_),
    .A1(\cpuregs[3][4] ),
    .S(_13931_),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_1 _17325_ (.A0(_13921_),
    .A1(\cpuregs[3][3] ),
    .S(_13931_),
    .X(_03410_));
 sky130_fd_sc_hd__mux2_1 _17326_ (.A0(_13922_),
    .A1(\cpuregs[3][2] ),
    .S(_13931_),
    .X(_03409_));
 sky130_fd_sc_hd__mux2_1 _17327_ (.A0(_13923_),
    .A1(\cpuregs[3][1] ),
    .S(_13926_),
    .X(_03408_));
 sky130_fd_sc_hd__mux2_1 _17328_ (.A0(_13924_),
    .A1(\cpuregs[3][0] ),
    .S(_13926_),
    .X(_03407_));
 sky130_fd_sc_hd__and2_1 _17329_ (.A(_13786_),
    .B(_13738_),
    .X(_13932_));
 sky130_fd_sc_hd__buf_6 _17330_ (.A(_13932_),
    .X(_13933_));
 sky130_fd_sc_hd__clkbuf_4 _17331_ (.A(_13933_),
    .X(_13934_));
 sky130_fd_sc_hd__mux2_1 _17332_ (.A0(\cpuregs[1][31] ),
    .A1(\cpuregs_wrdata[31] ),
    .S(_13934_),
    .X(_03406_));
 sky130_fd_sc_hd__mux2_1 _17333_ (.A0(\cpuregs[1][30] ),
    .A1(\cpuregs_wrdata[30] ),
    .S(_13934_),
    .X(_03405_));
 sky130_fd_sc_hd__mux2_1 _17334_ (.A0(\cpuregs[1][29] ),
    .A1(\cpuregs_wrdata[29] ),
    .S(_13934_),
    .X(_03404_));
 sky130_fd_sc_hd__mux2_1 _17335_ (.A0(\cpuregs[1][28] ),
    .A1(\cpuregs_wrdata[28] ),
    .S(_13934_),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _17336_ (.A0(\cpuregs[1][27] ),
    .A1(\cpuregs_wrdata[27] ),
    .S(_13934_),
    .X(_03402_));
 sky130_fd_sc_hd__mux2_1 _17337_ (.A0(\cpuregs[1][26] ),
    .A1(\cpuregs_wrdata[26] ),
    .S(_13934_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_4 _17338_ (.A(_13933_),
    .X(_13935_));
 sky130_fd_sc_hd__mux2_1 _17339_ (.A0(\cpuregs[1][25] ),
    .A1(\cpuregs_wrdata[25] ),
    .S(_13935_),
    .X(_03400_));
 sky130_fd_sc_hd__mux2_1 _17340_ (.A0(\cpuregs[1][24] ),
    .A1(\cpuregs_wrdata[24] ),
    .S(_13935_),
    .X(_03399_));
 sky130_fd_sc_hd__mux2_1 _17341_ (.A0(\cpuregs[1][23] ),
    .A1(\cpuregs_wrdata[23] ),
    .S(_13935_),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_1 _17342_ (.A0(\cpuregs[1][22] ),
    .A1(\cpuregs_wrdata[22] ),
    .S(_13935_),
    .X(_03397_));
 sky130_fd_sc_hd__mux2_1 _17343_ (.A0(\cpuregs[1][21] ),
    .A1(\cpuregs_wrdata[21] ),
    .S(_13935_),
    .X(_03396_));
 sky130_fd_sc_hd__mux2_1 _17344_ (.A0(\cpuregs[1][20] ),
    .A1(\cpuregs_wrdata[20] ),
    .S(_13935_),
    .X(_03395_));
 sky130_fd_sc_hd__clkbuf_4 _17345_ (.A(_13933_),
    .X(_13936_));
 sky130_fd_sc_hd__mux2_1 _17346_ (.A0(\cpuregs[1][19] ),
    .A1(\cpuregs_wrdata[19] ),
    .S(_13936_),
    .X(_03394_));
 sky130_fd_sc_hd__mux2_1 _17347_ (.A0(\cpuregs[1][18] ),
    .A1(\cpuregs_wrdata[18] ),
    .S(_13936_),
    .X(_03393_));
 sky130_fd_sc_hd__mux2_1 _17348_ (.A0(\cpuregs[1][17] ),
    .A1(\cpuregs_wrdata[17] ),
    .S(_13936_),
    .X(_03392_));
 sky130_fd_sc_hd__mux2_1 _17349_ (.A0(\cpuregs[1][16] ),
    .A1(\cpuregs_wrdata[16] ),
    .S(_13936_),
    .X(_03391_));
 sky130_fd_sc_hd__mux2_1 _17350_ (.A0(\cpuregs[1][15] ),
    .A1(\cpuregs_wrdata[15] ),
    .S(_13936_),
    .X(_03390_));
 sky130_fd_sc_hd__mux2_1 _17351_ (.A0(\cpuregs[1][14] ),
    .A1(\cpuregs_wrdata[14] ),
    .S(_13936_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_4 _17352_ (.A(_13933_),
    .X(_13937_));
 sky130_fd_sc_hd__mux2_1 _17353_ (.A0(\cpuregs[1][13] ),
    .A1(\cpuregs_wrdata[13] ),
    .S(_13937_),
    .X(_03388_));
 sky130_fd_sc_hd__mux2_1 _17354_ (.A0(\cpuregs[1][12] ),
    .A1(\cpuregs_wrdata[12] ),
    .S(_13937_),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _17355_ (.A0(\cpuregs[1][11] ),
    .A1(\cpuregs_wrdata[11] ),
    .S(_13937_),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_1 _17356_ (.A0(\cpuregs[1][10] ),
    .A1(\cpuregs_wrdata[10] ),
    .S(_13937_),
    .X(_03385_));
 sky130_fd_sc_hd__mux2_1 _17357_ (.A0(\cpuregs[1][9] ),
    .A1(\cpuregs_wrdata[9] ),
    .S(_13937_),
    .X(_03384_));
 sky130_fd_sc_hd__mux2_1 _17358_ (.A0(\cpuregs[1][8] ),
    .A1(\cpuregs_wrdata[8] ),
    .S(_13937_),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_4 _17359_ (.A(_13932_),
    .X(_13938_));
 sky130_fd_sc_hd__mux2_1 _17360_ (.A0(\cpuregs[1][7] ),
    .A1(\cpuregs_wrdata[7] ),
    .S(_13938_),
    .X(_03382_));
 sky130_fd_sc_hd__mux2_1 _17361_ (.A0(\cpuregs[1][6] ),
    .A1(\cpuregs_wrdata[6] ),
    .S(_13938_),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_1 _17362_ (.A0(\cpuregs[1][5] ),
    .A1(\cpuregs_wrdata[5] ),
    .S(_13938_),
    .X(_03380_));
 sky130_fd_sc_hd__mux2_1 _17363_ (.A0(\cpuregs[1][4] ),
    .A1(\cpuregs_wrdata[4] ),
    .S(_13938_),
    .X(_03379_));
 sky130_fd_sc_hd__mux2_1 _17364_ (.A0(\cpuregs[1][3] ),
    .A1(\cpuregs_wrdata[3] ),
    .S(_13938_),
    .X(_03378_));
 sky130_fd_sc_hd__mux2_1 _17365_ (.A0(\cpuregs[1][2] ),
    .A1(\cpuregs_wrdata[2] ),
    .S(_13938_),
    .X(_03377_));
 sky130_fd_sc_hd__mux2_1 _17366_ (.A0(\cpuregs[1][1] ),
    .A1(\cpuregs_wrdata[1] ),
    .S(_13933_),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_1 _17367_ (.A0(\cpuregs[1][0] ),
    .A1(\cpuregs_wrdata[0] ),
    .S(_13933_),
    .X(_03375_));
 sky130_fd_sc_hd__nand3b_2 _17368_ (.A_N(_13742_),
    .B(_13739_),
    .C(_13878_),
    .Y(_13939_));
 sky130_fd_sc_hd__buf_6 _17369_ (.A(_13939_),
    .X(_13940_));
 sky130_fd_sc_hd__clkbuf_4 _17370_ (.A(_13940_),
    .X(_13941_));
 sky130_fd_sc_hd__mux2_1 _17371_ (.A0(_13886_),
    .A1(\cpuregs[12][31] ),
    .S(_13941_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _17372_ (.A0(_13890_),
    .A1(\cpuregs[12][30] ),
    .S(_13941_),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_1 _17373_ (.A0(_13891_),
    .A1(\cpuregs[12][29] ),
    .S(_13941_),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_1 _17374_ (.A0(_13892_),
    .A1(\cpuregs[12][28] ),
    .S(_13941_),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_1 _17375_ (.A0(_13893_),
    .A1(\cpuregs[12][27] ),
    .S(_13941_),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_1 _17376_ (.A0(_13894_),
    .A1(\cpuregs[12][26] ),
    .S(_13941_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_4 _17377_ (.A(_13940_),
    .X(_13942_));
 sky130_fd_sc_hd__mux2_1 _17378_ (.A0(_13895_),
    .A1(\cpuregs[12][25] ),
    .S(_13942_),
    .X(_03368_));
 sky130_fd_sc_hd__mux2_1 _17379_ (.A0(_13897_),
    .A1(\cpuregs[12][24] ),
    .S(_13942_),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_1 _17380_ (.A0(_13898_),
    .A1(\cpuregs[12][23] ),
    .S(_13942_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_1 _17381_ (.A0(_13899_),
    .A1(\cpuregs[12][22] ),
    .S(_13942_),
    .X(_03365_));
 sky130_fd_sc_hd__mux2_1 _17382_ (.A0(_13900_),
    .A1(\cpuregs[12][21] ),
    .S(_13942_),
    .X(_03364_));
 sky130_fd_sc_hd__mux2_1 _17383_ (.A0(_13901_),
    .A1(\cpuregs[12][20] ),
    .S(_13942_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_4 _17384_ (.A(_13940_),
    .X(_13943_));
 sky130_fd_sc_hd__mux2_1 _17385_ (.A0(_13902_),
    .A1(\cpuregs[12][19] ),
    .S(_13943_),
    .X(_03362_));
 sky130_fd_sc_hd__mux2_1 _17386_ (.A0(_13904_),
    .A1(\cpuregs[12][18] ),
    .S(_13943_),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_1 _17387_ (.A0(_13905_),
    .A1(\cpuregs[12][17] ),
    .S(_13943_),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_1 _17388_ (.A0(_13906_),
    .A1(\cpuregs[12][16] ),
    .S(_13943_),
    .X(_03359_));
 sky130_fd_sc_hd__mux2_1 _17389_ (.A0(_13907_),
    .A1(\cpuregs[12][15] ),
    .S(_13943_),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_1 _17390_ (.A0(_13908_),
    .A1(\cpuregs[12][14] ),
    .S(_13943_),
    .X(_03357_));
 sky130_fd_sc_hd__buf_4 _17391_ (.A(_13940_),
    .X(_13944_));
 sky130_fd_sc_hd__mux2_1 _17392_ (.A0(_13909_),
    .A1(\cpuregs[12][13] ),
    .S(_13944_),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_1 _17393_ (.A0(_13911_),
    .A1(\cpuregs[12][12] ),
    .S(_13944_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _17394_ (.A0(_13912_),
    .A1(\cpuregs[12][11] ),
    .S(_13944_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_1 _17395_ (.A0(_13913_),
    .A1(\cpuregs[12][10] ),
    .S(_13944_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_1 _17396_ (.A0(_13914_),
    .A1(\cpuregs[12][9] ),
    .S(_13944_),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_1 _17397_ (.A0(_13915_),
    .A1(\cpuregs[12][8] ),
    .S(_13944_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_4 _17398_ (.A(_13939_),
    .X(_13945_));
 sky130_fd_sc_hd__mux2_1 _17399_ (.A0(_13916_),
    .A1(\cpuregs[12][7] ),
    .S(_13945_),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_1 _17400_ (.A0(_13918_),
    .A1(\cpuregs[12][6] ),
    .S(_13945_),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_1 _17401_ (.A0(_13919_),
    .A1(\cpuregs[12][5] ),
    .S(_13945_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _17402_ (.A0(_13920_),
    .A1(\cpuregs[12][4] ),
    .S(_13945_),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_1 _17403_ (.A0(_13921_),
    .A1(\cpuregs[12][3] ),
    .S(_13945_),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_1 _17404_ (.A0(_13922_),
    .A1(\cpuregs[12][2] ),
    .S(_13945_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _17405_ (.A0(_13923_),
    .A1(\cpuregs[12][1] ),
    .S(_13940_),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_1 _17406_ (.A0(_13924_),
    .A1(\cpuregs[12][0] ),
    .S(_13940_),
    .X(_03343_));
 sky130_fd_sc_hd__nor3_1 _17407_ (.A(\latched_rd[0] ),
    .B(\latched_rd[1] ),
    .C(_13742_),
    .Y(_13946_));
 sky130_fd_sc_hd__or3b_4 _17408_ (.A(_13745_),
    .B(_13744_),
    .C_N(_13946_),
    .X(_13947_));
 sky130_fd_sc_hd__buf_6 _17409_ (.A(_13947_),
    .X(_13948_));
 sky130_fd_sc_hd__clkbuf_4 _17410_ (.A(_13948_),
    .X(_13949_));
 sky130_fd_sc_hd__mux2_1 _17411_ (.A0(_13886_),
    .A1(\cpuregs[16][31] ),
    .S(_13949_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_1 _17412_ (.A0(_13890_),
    .A1(\cpuregs[16][30] ),
    .S(_13949_),
    .X(_03341_));
 sky130_fd_sc_hd__mux2_1 _17413_ (.A0(_13891_),
    .A1(\cpuregs[16][29] ),
    .S(_13949_),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_1 _17414_ (.A0(_13892_),
    .A1(\cpuregs[16][28] ),
    .S(_13949_),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _17415_ (.A0(_13893_),
    .A1(\cpuregs[16][27] ),
    .S(_13949_),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_1 _17416_ (.A0(_13894_),
    .A1(\cpuregs[16][26] ),
    .S(_13949_),
    .X(_03337_));
 sky130_fd_sc_hd__clkbuf_4 _17417_ (.A(_13948_),
    .X(_13950_));
 sky130_fd_sc_hd__mux2_1 _17418_ (.A0(_13895_),
    .A1(\cpuregs[16][25] ),
    .S(_13950_),
    .X(_03336_));
 sky130_fd_sc_hd__mux2_1 _17419_ (.A0(_13897_),
    .A1(\cpuregs[16][24] ),
    .S(_13950_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _17420_ (.A0(_13898_),
    .A1(\cpuregs[16][23] ),
    .S(_13950_),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_1 _17421_ (.A0(_13899_),
    .A1(\cpuregs[16][22] ),
    .S(_13950_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _17422_ (.A0(_13900_),
    .A1(\cpuregs[16][21] ),
    .S(_13950_),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_1 _17423_ (.A0(_13901_),
    .A1(\cpuregs[16][20] ),
    .S(_13950_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_4 _17424_ (.A(_13948_),
    .X(_13951_));
 sky130_fd_sc_hd__mux2_1 _17425_ (.A0(_13902_),
    .A1(\cpuregs[16][19] ),
    .S(_13951_),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_1 _17426_ (.A0(_13904_),
    .A1(\cpuregs[16][18] ),
    .S(_13951_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_1 _17427_ (.A0(_13905_),
    .A1(\cpuregs[16][17] ),
    .S(_13951_),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_1 _17428_ (.A0(_13906_),
    .A1(\cpuregs[16][16] ),
    .S(_13951_),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_1 _17429_ (.A0(_13907_),
    .A1(\cpuregs[16][15] ),
    .S(_13951_),
    .X(_03326_));
 sky130_fd_sc_hd__mux2_1 _17430_ (.A0(_13908_),
    .A1(\cpuregs[16][14] ),
    .S(_13951_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_4 _17431_ (.A(_13948_),
    .X(_13952_));
 sky130_fd_sc_hd__mux2_1 _17432_ (.A0(_13909_),
    .A1(\cpuregs[16][13] ),
    .S(_13952_),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_1 _17433_ (.A0(_13911_),
    .A1(\cpuregs[16][12] ),
    .S(_13952_),
    .X(_03323_));
 sky130_fd_sc_hd__mux2_1 _17434_ (.A0(_13912_),
    .A1(\cpuregs[16][11] ),
    .S(_13952_),
    .X(_03322_));
 sky130_fd_sc_hd__mux2_1 _17435_ (.A0(_13913_),
    .A1(\cpuregs[16][10] ),
    .S(_13952_),
    .X(_03321_));
 sky130_fd_sc_hd__mux2_1 _17436_ (.A0(_13914_),
    .A1(\cpuregs[16][9] ),
    .S(_13952_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _17437_ (.A0(_13915_),
    .A1(\cpuregs[16][8] ),
    .S(_13952_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_4 _17438_ (.A(_13947_),
    .X(_13953_));
 sky130_fd_sc_hd__mux2_1 _17439_ (.A0(_13916_),
    .A1(\cpuregs[16][7] ),
    .S(_13953_),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_1 _17440_ (.A0(_13918_),
    .A1(\cpuregs[16][6] ),
    .S(_13953_),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_1 _17441_ (.A0(_13919_),
    .A1(\cpuregs[16][5] ),
    .S(_13953_),
    .X(_03316_));
 sky130_fd_sc_hd__mux2_1 _17442_ (.A0(_13920_),
    .A1(\cpuregs[16][4] ),
    .S(_13953_),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_1 _17443_ (.A0(_13921_),
    .A1(\cpuregs[16][3] ),
    .S(_13953_),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_1 _17444_ (.A0(_13922_),
    .A1(\cpuregs[16][2] ),
    .S(_13953_),
    .X(_03313_));
 sky130_fd_sc_hd__mux2_1 _17445_ (.A0(_13923_),
    .A1(\cpuregs[16][1] ),
    .S(_13948_),
    .X(_03312_));
 sky130_fd_sc_hd__mux2_1 _17446_ (.A0(_13924_),
    .A1(\cpuregs[16][0] ),
    .S(_13948_),
    .X(_03311_));
 sky130_fd_sc_hd__nand2_1 _17447_ (.A(_13786_),
    .B(_13849_),
    .Y(_13954_));
 sky130_fd_sc_hd__buf_6 _17448_ (.A(_13954_),
    .X(_13955_));
 sky130_fd_sc_hd__clkbuf_4 _17449_ (.A(_13955_),
    .X(_13956_));
 sky130_fd_sc_hd__mux2_1 _17450_ (.A0(_13886_),
    .A1(\cpuregs[17][31] ),
    .S(_13956_),
    .X(_03310_));
 sky130_fd_sc_hd__mux2_1 _17451_ (.A0(_13890_),
    .A1(\cpuregs[17][30] ),
    .S(_13956_),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_1 _17452_ (.A0(_13891_),
    .A1(\cpuregs[17][29] ),
    .S(_13956_),
    .X(_03308_));
 sky130_fd_sc_hd__mux2_1 _17453_ (.A0(_13892_),
    .A1(\cpuregs[17][28] ),
    .S(_13956_),
    .X(_03307_));
 sky130_fd_sc_hd__mux2_1 _17454_ (.A0(_13893_),
    .A1(\cpuregs[17][27] ),
    .S(_13956_),
    .X(_03306_));
 sky130_fd_sc_hd__mux2_1 _17455_ (.A0(_13894_),
    .A1(\cpuregs[17][26] ),
    .S(_13956_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_4 _17456_ (.A(_13955_),
    .X(_13957_));
 sky130_fd_sc_hd__mux2_1 _17457_ (.A0(_13895_),
    .A1(\cpuregs[17][25] ),
    .S(_13957_),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_1 _17458_ (.A0(_13897_),
    .A1(\cpuregs[17][24] ),
    .S(_13957_),
    .X(_03303_));
 sky130_fd_sc_hd__mux2_1 _17459_ (.A0(_13898_),
    .A1(\cpuregs[17][23] ),
    .S(_13957_),
    .X(_03302_));
 sky130_fd_sc_hd__mux2_1 _17460_ (.A0(_13899_),
    .A1(\cpuregs[17][22] ),
    .S(_13957_),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_1 _17461_ (.A0(_13900_),
    .A1(\cpuregs[17][21] ),
    .S(_13957_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_1 _17462_ (.A0(_13901_),
    .A1(\cpuregs[17][20] ),
    .S(_13957_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_4 _17463_ (.A(_13955_),
    .X(_13958_));
 sky130_fd_sc_hd__mux2_1 _17464_ (.A0(_13902_),
    .A1(\cpuregs[17][19] ),
    .S(_13958_),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_1 _17465_ (.A0(_13904_),
    .A1(\cpuregs[17][18] ),
    .S(_13958_),
    .X(_03297_));
 sky130_fd_sc_hd__mux2_1 _17466_ (.A0(_13905_),
    .A1(\cpuregs[17][17] ),
    .S(_13958_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _17467_ (.A0(_13906_),
    .A1(\cpuregs[17][16] ),
    .S(_13958_),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_1 _17468_ (.A0(_13907_),
    .A1(\cpuregs[17][15] ),
    .S(_13958_),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_1 _17469_ (.A0(_13908_),
    .A1(\cpuregs[17][14] ),
    .S(_13958_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_4 _17470_ (.A(_13955_),
    .X(_13959_));
 sky130_fd_sc_hd__mux2_1 _17471_ (.A0(_13909_),
    .A1(\cpuregs[17][13] ),
    .S(_13959_),
    .X(_03292_));
 sky130_fd_sc_hd__mux2_1 _17472_ (.A0(_13911_),
    .A1(\cpuregs[17][12] ),
    .S(_13959_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _17473_ (.A0(_13912_),
    .A1(\cpuregs[17][11] ),
    .S(_13959_),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _17474_ (.A0(_13913_),
    .A1(\cpuregs[17][10] ),
    .S(_13959_),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_1 _17475_ (.A0(_13914_),
    .A1(\cpuregs[17][9] ),
    .S(_13959_),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_1 _17476_ (.A0(_13915_),
    .A1(\cpuregs[17][8] ),
    .S(_13959_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_4 _17477_ (.A(_13954_),
    .X(_13960_));
 sky130_fd_sc_hd__mux2_1 _17478_ (.A0(_13916_),
    .A1(\cpuregs[17][7] ),
    .S(_13960_),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_1 _17479_ (.A0(_13918_),
    .A1(\cpuregs[17][6] ),
    .S(_13960_),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_1 _17480_ (.A0(_13919_),
    .A1(\cpuregs[17][5] ),
    .S(_13960_),
    .X(_03284_));
 sky130_fd_sc_hd__mux2_1 _17481_ (.A0(_13920_),
    .A1(\cpuregs[17][4] ),
    .S(_13960_),
    .X(_03283_));
 sky130_fd_sc_hd__mux2_1 _17482_ (.A0(_13921_),
    .A1(\cpuregs[17][3] ),
    .S(_13960_),
    .X(_03282_));
 sky130_fd_sc_hd__mux2_1 _17483_ (.A0(_13922_),
    .A1(\cpuregs[17][2] ),
    .S(_13960_),
    .X(_03281_));
 sky130_fd_sc_hd__mux2_1 _17484_ (.A0(_13923_),
    .A1(\cpuregs[17][1] ),
    .S(_13955_),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_1 _17485_ (.A0(_13924_),
    .A1(\cpuregs[17][0] ),
    .S(_13955_),
    .X(_03279_));
 sky130_fd_sc_hd__buf_4 _17486_ (.A(\pcpi_mul.rs2[31] ),
    .X(_13961_));
 sky130_fd_sc_hd__clkbuf_4 _17487_ (.A(_13961_),
    .X(_13962_));
 sky130_fd_sc_hd__buf_4 _17488_ (.A(_13962_),
    .X(_13963_));
 sky130_vsdinv _17489_ (.A(_12796_),
    .Y(_13964_));
 sky130_fd_sc_hd__and2_1 _17490_ (.A(_12807_),
    .B(_12808_),
    .X(_13965_));
 sky130_fd_sc_hd__a21o_1 _17491_ (.A1(_13963_),
    .A2(_13964_),
    .B1(_13965_),
    .X(_03278_));
 sky130_fd_sc_hd__clkinv_4 _17492_ (.A(\pcpi_mul.rs2[30] ),
    .Y(_13966_));
 sky130_fd_sc_hd__clkbuf_8 _17493_ (.A(_13966_),
    .X(_13967_));
 sky130_fd_sc_hd__buf_6 _17494_ (.A(_13967_),
    .X(_13968_));
 sky130_fd_sc_hd__buf_6 _17495_ (.A(_13968_),
    .X(_13969_));
 sky130_fd_sc_hd__nand2_1 _17496_ (.A(_12794_),
    .B(_13797_),
    .Y(_13970_));
 sky130_fd_sc_hd__o21ai_1 _17497_ (.A1(_13969_),
    .A2(_03728_),
    .B1(_13970_),
    .Y(_03277_));
 sky130_fd_sc_hd__buf_4 _17498_ (.A(\pcpi_mul.rs2[29] ),
    .X(_13971_));
 sky130_fd_sc_hd__buf_4 _17499_ (.A(_13971_),
    .X(_13972_));
 sky130_fd_sc_hd__buf_4 _17500_ (.A(_13972_),
    .X(_13973_));
 sky130_fd_sc_hd__buf_6 _17501_ (.A(_13973_),
    .X(_13974_));
 sky130_fd_sc_hd__and2_1 _17502_ (.A(_12807_),
    .B(_13798_),
    .X(_13975_));
 sky130_fd_sc_hd__a21o_1 _17503_ (.A1(_13974_),
    .A2(_13964_),
    .B1(_13975_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_2 _17504_ (.A(\pcpi_mul.rs2[28] ),
    .X(_13976_));
 sky130_fd_sc_hd__buf_2 _17505_ (.A(_13976_),
    .X(_13977_));
 sky130_fd_sc_hd__buf_6 _17506_ (.A(_13977_),
    .X(_13978_));
 sky130_fd_sc_hd__clkbuf_4 _17507_ (.A(_13978_),
    .X(_13979_));
 sky130_fd_sc_hd__buf_4 _17508_ (.A(_13979_),
    .X(_13980_));
 sky130_fd_sc_hd__and2_1 _17509_ (.A(_12807_),
    .B(_13799_),
    .X(_13981_));
 sky130_fd_sc_hd__a21o_1 _17510_ (.A1(_13980_),
    .A2(_13964_),
    .B1(_13981_),
    .X(_03275_));
 sky130_vsdinv _17511_ (.A(\pcpi_mul.rs2[27] ),
    .Y(_13982_));
 sky130_fd_sc_hd__nand2_1 _17512_ (.A(_12794_),
    .B(_13800_),
    .Y(_13983_));
 sky130_fd_sc_hd__o21ai_1 _17513_ (.A1(_13982_),
    .A2(_03728_),
    .B1(_13983_),
    .Y(_03274_));
 sky130_vsdinv _17514_ (.A(\pcpi_mul.rs2[26] ),
    .Y(_13984_));
 sky130_fd_sc_hd__buf_4 _17515_ (.A(_13984_),
    .X(_13985_));
 sky130_fd_sc_hd__buf_4 _17516_ (.A(_13985_),
    .X(_13986_));
 sky130_fd_sc_hd__nand2_1 _17517_ (.A(_12794_),
    .B(_13801_),
    .Y(_13987_));
 sky130_fd_sc_hd__o21ai_1 _17518_ (.A1(_13986_),
    .A2(_03728_),
    .B1(_13987_),
    .Y(_03273_));
 sky130_vsdinv _17519_ (.A(\pcpi_mul.rs2[25] ),
    .Y(_13988_));
 sky130_fd_sc_hd__buf_2 _17520_ (.A(_13988_),
    .X(_13989_));
 sky130_fd_sc_hd__buf_2 _17521_ (.A(_13989_),
    .X(_13990_));
 sky130_fd_sc_hd__buf_6 _17522_ (.A(_13990_),
    .X(_13991_));
 sky130_fd_sc_hd__nand2_1 _17523_ (.A(_12794_),
    .B(_13804_),
    .Y(_13992_));
 sky130_fd_sc_hd__o21ai_1 _17524_ (.A1(_13991_),
    .A2(_03728_),
    .B1(_13992_),
    .Y(_03272_));
 sky130_fd_sc_hd__clkinv_4 _17525_ (.A(\pcpi_mul.rs2[24] ),
    .Y(_13993_));
 sky130_fd_sc_hd__buf_4 _17526_ (.A(_12796_),
    .X(_13994_));
 sky130_fd_sc_hd__buf_2 _17527_ (.A(_12793_),
    .X(_13995_));
 sky130_fd_sc_hd__nand2_4 _17528_ (.A(_13995_),
    .B(_13805_),
    .Y(_13996_));
 sky130_fd_sc_hd__o21ai_1 _17529_ (.A1(_13993_),
    .A2(_13994_),
    .B1(_13996_),
    .Y(_03271_));
 sky130_fd_sc_hd__buf_2 _17530_ (.A(\pcpi_mul.rs2[23] ),
    .X(_13997_));
 sky130_fd_sc_hd__clkbuf_4 _17531_ (.A(_13997_),
    .X(_13998_));
 sky130_vsdinv _17532_ (.A(_13998_),
    .Y(_13999_));
 sky130_fd_sc_hd__nand2_2 _17533_ (.A(_13995_),
    .B(_13806_),
    .Y(_14000_));
 sky130_fd_sc_hd__o21ai_1 _17534_ (.A1(_13999_),
    .A2(_13994_),
    .B1(_14000_),
    .Y(_03270_));
 sky130_fd_sc_hd__buf_4 _17535_ (.A(\pcpi_mul.rs2[22] ),
    .X(_14001_));
 sky130_vsdinv _17536_ (.A(_14001_),
    .Y(_14002_));
 sky130_fd_sc_hd__nand2_2 _17537_ (.A(_13995_),
    .B(_13807_),
    .Y(_14003_));
 sky130_fd_sc_hd__o21ai_1 _17538_ (.A1(_14002_),
    .A2(_13994_),
    .B1(_14003_),
    .Y(_03269_));
 sky130_vsdinv _17539_ (.A(\pcpi_mul.rs2[21] ),
    .Y(_14004_));
 sky130_fd_sc_hd__buf_2 _17540_ (.A(_14004_),
    .X(_14005_));
 sky130_fd_sc_hd__clkbuf_8 _17541_ (.A(_14005_),
    .X(_14006_));
 sky130_fd_sc_hd__nand2_1 _17542_ (.A(_13995_),
    .B(_13808_),
    .Y(_14007_));
 sky130_fd_sc_hd__o21ai_1 _17543_ (.A1(_14006_),
    .A2(_13994_),
    .B1(_14007_),
    .Y(_03268_));
 sky130_fd_sc_hd__buf_2 _17544_ (.A(\pcpi_mul.rs2[20] ),
    .X(_14008_));
 sky130_fd_sc_hd__buf_4 _17545_ (.A(_14008_),
    .X(_14009_));
 sky130_fd_sc_hd__buf_4 _17546_ (.A(_14009_),
    .X(_14010_));
 sky130_vsdinv _17547_ (.A(_14010_),
    .Y(_14011_));
 sky130_fd_sc_hd__nand2_2 _17548_ (.A(_13995_),
    .B(_13809_),
    .Y(_14012_));
 sky130_fd_sc_hd__o21ai_2 _17549_ (.A1(_14011_),
    .A2(_13994_),
    .B1(_14012_),
    .Y(_03267_));
 sky130_fd_sc_hd__buf_2 _17550_ (.A(\pcpi_mul.rs2[19] ),
    .X(_14013_));
 sky130_fd_sc_hd__clkbuf_4 _17551_ (.A(_14013_),
    .X(_14014_));
 sky130_fd_sc_hd__buf_4 _17552_ (.A(_14014_),
    .X(_14015_));
 sky130_vsdinv _17553_ (.A(_14015_),
    .Y(_14016_));
 sky130_fd_sc_hd__nand2_2 _17554_ (.A(_13995_),
    .B(_13811_),
    .Y(_14017_));
 sky130_fd_sc_hd__o21ai_2 _17555_ (.A1(_14016_),
    .A2(_13994_),
    .B1(_14017_),
    .Y(_03266_));
 sky130_vsdinv _17556_ (.A(\pcpi_mul.rs2[18] ),
    .Y(_14018_));
 sky130_fd_sc_hd__clkbuf_4 _17557_ (.A(_12796_),
    .X(_14019_));
 sky130_fd_sc_hd__clkbuf_4 _17558_ (.A(_12793_),
    .X(_14020_));
 sky130_fd_sc_hd__nand2_4 _17559_ (.A(_14020_),
    .B(_13812_),
    .Y(_14021_));
 sky130_fd_sc_hd__o21ai_4 _17560_ (.A1(_14018_),
    .A2(_14019_),
    .B1(_14021_),
    .Y(_03265_));
 sky130_fd_sc_hd__clkbuf_2 _17561_ (.A(\pcpi_mul.rs2[17] ),
    .X(_14022_));
 sky130_fd_sc_hd__buf_2 _17562_ (.A(_14022_),
    .X(_14023_));
 sky130_vsdinv _17563_ (.A(_14023_),
    .Y(_14024_));
 sky130_fd_sc_hd__nand2_2 _17564_ (.A(_14020_),
    .B(_13813_),
    .Y(_14025_));
 sky130_fd_sc_hd__o21ai_2 _17565_ (.A1(_14024_),
    .A2(_14019_),
    .B1(_14025_),
    .Y(_03264_));
 sky130_fd_sc_hd__clkbuf_4 _17566_ (.A(\pcpi_mul.rs2[16] ),
    .X(_14026_));
 sky130_fd_sc_hd__clkbuf_4 _17567_ (.A(_14026_),
    .X(_14027_));
 sky130_vsdinv _17568_ (.A(_14027_),
    .Y(_14028_));
 sky130_fd_sc_hd__nand2_2 _17569_ (.A(_14020_),
    .B(_13814_),
    .Y(_14029_));
 sky130_fd_sc_hd__o21ai_1 _17570_ (.A1(_14028_),
    .A2(_14019_),
    .B1(_14029_),
    .Y(_03263_));
 sky130_vsdinv _17571_ (.A(\pcpi_mul.rs2[15] ),
    .Y(_14030_));
 sky130_fd_sc_hd__buf_2 _17572_ (.A(_14030_),
    .X(_14031_));
 sky130_fd_sc_hd__buf_4 _17573_ (.A(_14031_),
    .X(_14032_));
 sky130_fd_sc_hd__buf_6 _17574_ (.A(_14032_),
    .X(_14033_));
 sky130_fd_sc_hd__nand2_2 _17575_ (.A(_14020_),
    .B(_13815_),
    .Y(_14034_));
 sky130_fd_sc_hd__o21ai_2 _17576_ (.A1(_14033_),
    .A2(_14019_),
    .B1(_14034_),
    .Y(_03262_));
 sky130_fd_sc_hd__clkbuf_4 _17577_ (.A(\pcpi_mul.rs2[14] ),
    .X(_14035_));
 sky130_fd_sc_hd__buf_4 _17578_ (.A(_14035_),
    .X(_14036_));
 sky130_fd_sc_hd__buf_6 _17579_ (.A(_14036_),
    .X(_14037_));
 sky130_fd_sc_hd__buf_8 _17580_ (.A(_14037_),
    .X(_14038_));
 sky130_fd_sc_hd__and2_1 _17581_ (.A(_12807_),
    .B(_13816_),
    .X(_14039_));
 sky130_fd_sc_hd__a21o_1 _17582_ (.A1(_14038_),
    .A2(_13964_),
    .B1(_14039_),
    .X(_03261_));
 sky130_fd_sc_hd__clkbuf_4 _17583_ (.A(\pcpi_mul.rs2[13] ),
    .X(_14040_));
 sky130_fd_sc_hd__buf_4 _17584_ (.A(_14040_),
    .X(_14041_));
 sky130_fd_sc_hd__buf_4 _17585_ (.A(_14041_),
    .X(_14042_));
 sky130_fd_sc_hd__buf_8 _17586_ (.A(_14042_),
    .X(_14043_));
 sky130_fd_sc_hd__and2_1 _17587_ (.A(_12807_),
    .B(_13818_),
    .X(_14044_));
 sky130_fd_sc_hd__a21o_1 _17588_ (.A1(_14043_),
    .A2(_13964_),
    .B1(_14044_),
    .X(_03260_));
 sky130_vsdinv _17589_ (.A(\pcpi_mul.rs2[12] ),
    .Y(_14045_));
 sky130_fd_sc_hd__buf_4 _17590_ (.A(_14045_),
    .X(_14046_));
 sky130_fd_sc_hd__buf_4 _17591_ (.A(_14046_),
    .X(_14047_));
 sky130_fd_sc_hd__clkbuf_4 _17592_ (.A(_14047_),
    .X(_14048_));
 sky130_fd_sc_hd__nand2_2 _17593_ (.A(_14020_),
    .B(_13819_),
    .Y(_14049_));
 sky130_fd_sc_hd__o21ai_1 _17594_ (.A1(_14048_),
    .A2(_14019_),
    .B1(_14049_),
    .Y(_03259_));
 sky130_fd_sc_hd__buf_4 _17595_ (.A(\pcpi_mul.rs2[11] ),
    .X(_14050_));
 sky130_vsdinv _17596_ (.A(_14050_),
    .Y(_14051_));
 sky130_fd_sc_hd__nand2_2 _17597_ (.A(_14020_),
    .B(_13820_),
    .Y(_14052_));
 sky130_fd_sc_hd__o21ai_1 _17598_ (.A1(_14051_),
    .A2(_14019_),
    .B1(_14052_),
    .Y(_03258_));
 sky130_fd_sc_hd__clkbuf_4 _17599_ (.A(\pcpi_mul.rs2[10] ),
    .X(_14053_));
 sky130_vsdinv _17600_ (.A(_14053_),
    .Y(_14054_));
 sky130_fd_sc_hd__clkbuf_2 _17601_ (.A(_12796_),
    .X(_14055_));
 sky130_fd_sc_hd__buf_2 _17602_ (.A(_12793_),
    .X(_14056_));
 sky130_fd_sc_hd__nand2_2 _17603_ (.A(_14056_),
    .B(_13821_),
    .Y(_14057_));
 sky130_fd_sc_hd__o21ai_1 _17604_ (.A1(_14054_),
    .A2(_14055_),
    .B1(_14057_),
    .Y(_03257_));
 sky130_vsdinv _17605_ (.A(\pcpi_mul.rs2[9] ),
    .Y(_14058_));
 sky130_fd_sc_hd__clkbuf_4 _17606_ (.A(_14058_),
    .X(_14059_));
 sky130_fd_sc_hd__nand2_2 _17607_ (.A(_14056_),
    .B(_13822_),
    .Y(_14060_));
 sky130_fd_sc_hd__o21ai_1 _17608_ (.A1(_14059_),
    .A2(_14055_),
    .B1(_14060_),
    .Y(_03256_));
 sky130_fd_sc_hd__clkbuf_4 _17609_ (.A(\pcpi_mul.rs2[8] ),
    .X(_14061_));
 sky130_fd_sc_hd__buf_4 _17610_ (.A(_14061_),
    .X(_14062_));
 sky130_vsdinv _17611_ (.A(_14062_),
    .Y(_14063_));
 sky130_fd_sc_hd__nand2_1 _17612_ (.A(_14056_),
    .B(_13823_),
    .Y(_14064_));
 sky130_fd_sc_hd__o21ai_1 _17613_ (.A1(_14063_),
    .A2(_14055_),
    .B1(_14064_),
    .Y(_03255_));
 sky130_fd_sc_hd__clkbuf_4 _17614_ (.A(\pcpi_mul.rs2[7] ),
    .X(_14065_));
 sky130_fd_sc_hd__clkbuf_4 _17615_ (.A(_14065_),
    .X(_14066_));
 sky130_vsdinv _17616_ (.A(_14066_),
    .Y(_14067_));
 sky130_fd_sc_hd__nand2_1 _17617_ (.A(_14056_),
    .B(_13826_),
    .Y(_14068_));
 sky130_fd_sc_hd__o21ai_1 _17618_ (.A1(_14067_),
    .A2(_14055_),
    .B1(_14068_),
    .Y(_03254_));
 sky130_fd_sc_hd__inv_2 _17619_ (.A(\pcpi_mul.rs2[6] ),
    .Y(_14069_));
 sky130_fd_sc_hd__clkbuf_4 _17620_ (.A(_14069_),
    .X(_14070_));
 sky130_fd_sc_hd__buf_4 _17621_ (.A(_14070_),
    .X(_14071_));
 sky130_fd_sc_hd__nand2_2 _17622_ (.A(_14056_),
    .B(_13828_),
    .Y(_14072_));
 sky130_fd_sc_hd__o21ai_1 _17623_ (.A1(_14071_),
    .A2(_14055_),
    .B1(_14072_),
    .Y(_03253_));
 sky130_fd_sc_hd__clkbuf_4 _17624_ (.A(\pcpi_mul.rs2[5] ),
    .X(_14073_));
 sky130_vsdinv _17625_ (.A(_14073_),
    .Y(_14074_));
 sky130_fd_sc_hd__clkbuf_4 _17626_ (.A(_14074_),
    .X(_14075_));
 sky130_fd_sc_hd__nand2_2 _17627_ (.A(_14056_),
    .B(_13830_),
    .Y(_14076_));
 sky130_fd_sc_hd__o21ai_2 _17628_ (.A1(_14075_),
    .A2(_14055_),
    .B1(_14076_),
    .Y(_03252_));
 sky130_vsdinv _17629_ (.A(\pcpi_mul.rs2[4] ),
    .Y(_14077_));
 sky130_fd_sc_hd__clkbuf_4 _17630_ (.A(_12795_),
    .X(_14078_));
 sky130_fd_sc_hd__buf_2 _17631_ (.A(_14078_),
    .X(_14079_));
 sky130_fd_sc_hd__buf_2 _17632_ (.A(_12793_),
    .X(_14080_));
 sky130_fd_sc_hd__nand2_1 _17633_ (.A(_14080_),
    .B(_13832_),
    .Y(_14081_));
 sky130_fd_sc_hd__o21ai_1 _17634_ (.A1(_14077_),
    .A2(_14079_),
    .B1(_14081_),
    .Y(_03251_));
 sky130_fd_sc_hd__buf_2 _17635_ (.A(\pcpi_mul.rs2[3] ),
    .X(_14082_));
 sky130_fd_sc_hd__buf_2 _17636_ (.A(_14082_),
    .X(_14083_));
 sky130_fd_sc_hd__buf_4 _17637_ (.A(_14083_),
    .X(_14084_));
 sky130_fd_sc_hd__inv_4 _17638_ (.A(_14084_),
    .Y(_14085_));
 sky130_fd_sc_hd__buf_6 _17639_ (.A(_14085_),
    .X(_14086_));
 sky130_fd_sc_hd__buf_6 _17640_ (.A(_14086_),
    .X(_14087_));
 sky130_fd_sc_hd__buf_6 _17641_ (.A(_14087_),
    .X(_14088_));
 sky130_fd_sc_hd__nand2_1 _17642_ (.A(_14080_),
    .B(_13834_),
    .Y(_14089_));
 sky130_fd_sc_hd__o21ai_1 _17643_ (.A1(_14088_),
    .A2(_14079_),
    .B1(_14089_),
    .Y(_03250_));
 sky130_fd_sc_hd__clkbuf_4 _17644_ (.A(\pcpi_mul.rs2[2] ),
    .X(_14090_));
 sky130_vsdinv _17645_ (.A(_14090_),
    .Y(_14091_));
 sky130_fd_sc_hd__nand2_1 _17646_ (.A(_14080_),
    .B(_13836_),
    .Y(_14092_));
 sky130_fd_sc_hd__o21ai_1 _17647_ (.A1(_14091_),
    .A2(_14079_),
    .B1(_14092_),
    .Y(_03249_));
 sky130_fd_sc_hd__clkbuf_4 _17648_ (.A(\pcpi_mul.rs2[1] ),
    .X(_14093_));
 sky130_vsdinv _17649_ (.A(_14093_),
    .Y(_14094_));
 sky130_fd_sc_hd__nand2_1 _17650_ (.A(_14080_),
    .B(_13838_),
    .Y(_14095_));
 sky130_fd_sc_hd__o21ai_1 _17651_ (.A1(_14094_),
    .A2(_14079_),
    .B1(_14095_),
    .Y(_03248_));
 sky130_vsdinv _17652_ (.A(\pcpi_mul.rs2[0] ),
    .Y(_14096_));
 sky130_fd_sc_hd__clkbuf_4 _17653_ (.A(_14096_),
    .X(_14097_));
 sky130_fd_sc_hd__buf_6 _17654_ (.A(_14097_),
    .X(_14098_));
 sky130_fd_sc_hd__nand2_1 _17655_ (.A(_14080_),
    .B(_13840_),
    .Y(_14099_));
 sky130_fd_sc_hd__o21ai_1 _17656_ (.A1(_14098_),
    .A2(_14079_),
    .B1(_14099_),
    .Y(_03247_));
 sky130_fd_sc_hd__mux2_1 _17657_ (.A0(net273),
    .A1(_02541_),
    .S(_12676_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _17658_ (.A0(net272),
    .A1(_02540_),
    .S(_12676_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_1 _17659_ (.A0(net271),
    .A1(_02539_),
    .S(_12675_),
    .X(_03244_));
 sky130_fd_sc_hd__mux2_1 _17660_ (.A0(net270),
    .A1(_02538_),
    .S(_12675_),
    .X(_03243_));
 sky130_fd_sc_hd__clkbuf_2 _17661_ (.A(_12680_),
    .X(_14100_));
 sky130_fd_sc_hd__and4b_1 _17662_ (.A_N(_12683_),
    .B(_14100_),
    .C(_12682_),
    .D(_12686_),
    .X(_14101_));
 sky130_fd_sc_hd__a32o_1 _17663_ (.A1(_14101_),
    .A2(_00329_),
    .A3(_00328_),
    .B1(_13019_),
    .B2(_12984_),
    .X(_03242_));
 sky130_vsdinv _17664_ (.A(_13047_),
    .Y(_14102_));
 sky130_fd_sc_hd__nand3_1 _17665_ (.A(_14101_),
    .B(_12684_),
    .C(_00328_),
    .Y(_14103_));
 sky130_fd_sc_hd__o21ai_1 _17666_ (.A1(_14102_),
    .A2(_15210_),
    .B1(_14103_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _17667_ (.A(_13786_),
    .B(_13878_),
    .Y(_14104_));
 sky130_fd_sc_hd__buf_6 _17668_ (.A(_14104_),
    .X(_14105_));
 sky130_fd_sc_hd__clkbuf_4 _17669_ (.A(_14105_),
    .X(_14106_));
 sky130_fd_sc_hd__mux2_1 _17670_ (.A0(_13886_),
    .A1(\cpuregs[13][31] ),
    .S(_14106_),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_1 _17671_ (.A0(_13890_),
    .A1(\cpuregs[13][30] ),
    .S(_14106_),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_1 _17672_ (.A0(_13891_),
    .A1(\cpuregs[13][29] ),
    .S(_14106_),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_1 _17673_ (.A0(_13892_),
    .A1(\cpuregs[13][28] ),
    .S(_14106_),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_1 _17674_ (.A0(_13893_),
    .A1(\cpuregs[13][27] ),
    .S(_14106_),
    .X(_03236_));
 sky130_fd_sc_hd__mux2_1 _17675_ (.A0(_13894_),
    .A1(\cpuregs[13][26] ),
    .S(_14106_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_4 _17676_ (.A(_14105_),
    .X(_14107_));
 sky130_fd_sc_hd__mux2_1 _17677_ (.A0(_13895_),
    .A1(\cpuregs[13][25] ),
    .S(_14107_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _17678_ (.A0(_13897_),
    .A1(\cpuregs[13][24] ),
    .S(_14107_),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_1 _17679_ (.A0(_13898_),
    .A1(\cpuregs[13][23] ),
    .S(_14107_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _17680_ (.A0(_13899_),
    .A1(\cpuregs[13][22] ),
    .S(_14107_),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_1 _17681_ (.A0(_13900_),
    .A1(\cpuregs[13][21] ),
    .S(_14107_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _17682_ (.A0(_13901_),
    .A1(\cpuregs[13][20] ),
    .S(_14107_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_4 _17683_ (.A(_14105_),
    .X(_14108_));
 sky130_fd_sc_hd__mux2_1 _17684_ (.A0(_13902_),
    .A1(\cpuregs[13][19] ),
    .S(_14108_),
    .X(_03228_));
 sky130_fd_sc_hd__mux2_1 _17685_ (.A0(_13904_),
    .A1(\cpuregs[13][18] ),
    .S(_14108_),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_1 _17686_ (.A0(_13905_),
    .A1(\cpuregs[13][17] ),
    .S(_14108_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_1 _17687_ (.A0(_13906_),
    .A1(\cpuregs[13][16] ),
    .S(_14108_),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_1 _17688_ (.A0(_13907_),
    .A1(\cpuregs[13][15] ),
    .S(_14108_),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_1 _17689_ (.A0(_13908_),
    .A1(\cpuregs[13][14] ),
    .S(_14108_),
    .X(_03223_));
 sky130_fd_sc_hd__buf_4 _17690_ (.A(_14105_),
    .X(_14109_));
 sky130_fd_sc_hd__mux2_1 _17691_ (.A0(_13909_),
    .A1(\cpuregs[13][13] ),
    .S(_14109_),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_1 _17692_ (.A0(_13911_),
    .A1(\cpuregs[13][12] ),
    .S(_14109_),
    .X(_03221_));
 sky130_fd_sc_hd__mux2_1 _17693_ (.A0(_13912_),
    .A1(\cpuregs[13][11] ),
    .S(_14109_),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_1 _17694_ (.A0(_13913_),
    .A1(\cpuregs[13][10] ),
    .S(_14109_),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_1 _17695_ (.A0(_13914_),
    .A1(\cpuregs[13][9] ),
    .S(_14109_),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_1 _17696_ (.A0(_13915_),
    .A1(\cpuregs[13][8] ),
    .S(_14109_),
    .X(_03217_));
 sky130_fd_sc_hd__buf_2 _17697_ (.A(_14104_),
    .X(_14110_));
 sky130_fd_sc_hd__mux2_1 _17698_ (.A0(_13916_),
    .A1(\cpuregs[13][7] ),
    .S(_14110_),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_1 _17699_ (.A0(_13918_),
    .A1(\cpuregs[13][6] ),
    .S(_14110_),
    .X(_03215_));
 sky130_fd_sc_hd__mux2_1 _17700_ (.A0(_13919_),
    .A1(\cpuregs[13][5] ),
    .S(_14110_),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_1 _17701_ (.A0(_13920_),
    .A1(\cpuregs[13][4] ),
    .S(_14110_),
    .X(_03213_));
 sky130_fd_sc_hd__mux2_1 _17702_ (.A0(_13921_),
    .A1(\cpuregs[13][3] ),
    .S(_14110_),
    .X(_03212_));
 sky130_fd_sc_hd__mux2_1 _17703_ (.A0(_13922_),
    .A1(\cpuregs[13][2] ),
    .S(_14110_),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_1 _17704_ (.A0(_13923_),
    .A1(\cpuregs[13][1] ),
    .S(_14105_),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_1 _17705_ (.A0(_13924_),
    .A1(\cpuregs[13][0] ),
    .S(_14105_),
    .X(_03209_));
 sky130_fd_sc_hd__buf_2 _17706_ (.A(is_sb_sh_sw),
    .X(_14111_));
 sky130_fd_sc_hd__clkbuf_4 _17707_ (.A(_14111_),
    .X(_14112_));
 sky130_fd_sc_hd__a32o_1 _17708_ (.A1(_14101_),
    .A2(_00329_),
    .A3(_12685_),
    .B1(_14112_),
    .B2(_12984_),
    .X(_03208_));
 sky130_fd_sc_hd__buf_2 _17709_ (.A(_13070_),
    .X(_14113_));
 sky130_fd_sc_hd__nor3b_2 _17710_ (.A(instr_jalr),
    .B(_13046_),
    .C_N(_13048_),
    .Y(_14114_));
 sky130_vsdinv _17711_ (.A(_13030_),
    .Y(_14115_));
 sky130_vsdinv _17712_ (.A(_13033_),
    .Y(_14116_));
 sky130_fd_sc_hd__a31o_1 _17713_ (.A1(_14115_),
    .A2(_00335_),
    .A3(_14116_),
    .B1(_14102_),
    .X(_14117_));
 sky130_fd_sc_hd__a2bb2oi_1 _17714_ (.A1_N(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2_N(_14113_),
    .B1(_14114_),
    .B2(_14117_),
    .Y(_03207_));
 sky130_fd_sc_hd__inv_2 _17715_ (.A(\mem_rdata_q[14] ),
    .Y(_00334_));
 sky130_fd_sc_hd__nor3_1 _17716_ (.A(_13014_),
    .B(_00334_),
    .C(_13017_),
    .Y(_14118_));
 sky130_fd_sc_hd__a31o_1 _17717_ (.A1(_12999_),
    .A2(_13000_),
    .A3(_12996_),
    .B1(_14118_),
    .X(_14119_));
 sky130_fd_sc_hd__and2b_1 _17718_ (.A_N(_12992_),
    .B(_12994_),
    .X(_14120_));
 sky130_fd_sc_hd__buf_2 _17719_ (.A(is_slli_srli_srai),
    .X(_14121_));
 sky130_fd_sc_hd__buf_2 _17720_ (.A(_13059_),
    .X(_14122_));
 sky130_fd_sc_hd__a32o_1 _17721_ (.A1(_14119_),
    .A2(_14120_),
    .A3(_13055_),
    .B1(_14121_),
    .B2(_14122_),
    .X(_03206_));
 sky130_fd_sc_hd__buf_2 _17722_ (.A(is_lb_lh_lw_lbu_lhu),
    .X(_14123_));
 sky130_fd_sc_hd__a32o_1 _17723_ (.A1(_14101_),
    .A2(_12684_),
    .A3(_12685_),
    .B1(_14123_),
    .B2(_12984_),
    .X(_03205_));
 sky130_fd_sc_hd__buf_6 _17724_ (.A(\decoded_imm_uj[20] ),
    .X(_14124_));
 sky130_fd_sc_hd__buf_4 _17725_ (.A(_14124_),
    .X(_14125_));
 sky130_fd_sc_hd__buf_6 _17726_ (.A(_14125_),
    .X(_14126_));
 sky130_fd_sc_hd__buf_2 _17727_ (.A(_14126_),
    .X(_14127_));
 sky130_fd_sc_hd__clkbuf_4 _17728_ (.A(_14100_),
    .X(_14128_));
 sky130_fd_sc_hd__mux2_1 _17729_ (.A0(_14127_),
    .A1(\mem_rdata_latched[31] ),
    .S(_14128_),
    .X(_03204_));
 sky130_fd_sc_hd__mux2_1 _17730_ (.A0(\decoded_imm_uj[19] ),
    .A1(\mem_rdata_latched[19] ),
    .S(_14128_),
    .X(_03203_));
 sky130_fd_sc_hd__mux2_1 _17731_ (.A0(\decoded_imm_uj[18] ),
    .A1(\mem_rdata_latched[18] ),
    .S(_14128_),
    .X(_03202_));
 sky130_fd_sc_hd__mux2_1 _17732_ (.A0(\decoded_imm_uj[17] ),
    .A1(\mem_rdata_latched[17] ),
    .S(_14128_),
    .X(_03201_));
 sky130_fd_sc_hd__mux2_1 _17733_ (.A0(\decoded_imm_uj[16] ),
    .A1(\mem_rdata_latched[16] ),
    .S(_14128_),
    .X(_03200_));
 sky130_fd_sc_hd__mux2_1 _17734_ (.A0(\decoded_imm_uj[15] ),
    .A1(\mem_rdata_latched[15] ),
    .S(_14128_),
    .X(_03199_));
 sky130_fd_sc_hd__buf_2 _17735_ (.A(_14100_),
    .X(_14129_));
 sky130_fd_sc_hd__mux2_1 _17736_ (.A0(\decoded_imm_uj[14] ),
    .A1(\mem_rdata_latched[14] ),
    .S(_14129_),
    .X(_03198_));
 sky130_fd_sc_hd__mux2_1 _17737_ (.A0(\decoded_imm_uj[13] ),
    .A1(\mem_rdata_latched[13] ),
    .S(_14129_),
    .X(_03197_));
 sky130_fd_sc_hd__mux2_1 _17738_ (.A0(\decoded_imm_uj[12] ),
    .A1(\mem_rdata_latched[12] ),
    .S(_14129_),
    .X(_03196_));
 sky130_fd_sc_hd__mux2_1 _17739_ (.A0(\decoded_imm_uj[11] ),
    .A1(\mem_rdata_latched[20] ),
    .S(_14129_),
    .X(_03195_));
 sky130_fd_sc_hd__mux2_1 _17740_ (.A0(\decoded_imm_uj[10] ),
    .A1(\mem_rdata_latched[30] ),
    .S(_14129_),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_1 _17741_ (.A0(\decoded_imm_uj[9] ),
    .A1(\mem_rdata_latched[29] ),
    .S(_14129_),
    .X(_03193_));
 sky130_fd_sc_hd__buf_2 _17742_ (.A(_14100_),
    .X(_14130_));
 sky130_fd_sc_hd__mux2_1 _17743_ (.A0(\decoded_imm_uj[8] ),
    .A1(\mem_rdata_latched[28] ),
    .S(_14130_),
    .X(_03192_));
 sky130_fd_sc_hd__mux2_1 _17744_ (.A0(\decoded_imm_uj[7] ),
    .A1(\mem_rdata_latched[27] ),
    .S(_14130_),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_1 _17745_ (.A0(\decoded_imm_uj[6] ),
    .A1(\mem_rdata_latched[26] ),
    .S(_14130_),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_1 _17746_ (.A0(\decoded_imm_uj[5] ),
    .A1(\mem_rdata_latched[25] ),
    .S(_14130_),
    .X(_03189_));
 sky130_fd_sc_hd__mux2_1 _17747_ (.A0(\decoded_imm_uj[4] ),
    .A1(\mem_rdata_latched[24] ),
    .S(_14130_),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_1 _17748_ (.A0(\decoded_imm_uj[3] ),
    .A1(\mem_rdata_latched[23] ),
    .S(_14130_),
    .X(_03187_));
 sky130_fd_sc_hd__clkbuf_4 _17749_ (.A(_14100_),
    .X(_14131_));
 sky130_fd_sc_hd__mux2_1 _17750_ (.A0(\decoded_imm_uj[2] ),
    .A1(\mem_rdata_latched[22] ),
    .S(_14131_),
    .X(_03186_));
 sky130_fd_sc_hd__mux2_1 _17751_ (.A0(\decoded_imm_uj[1] ),
    .A1(\mem_rdata_latched[21] ),
    .S(_14131_),
    .X(_03185_));
 sky130_vsdinv _17752_ (.A(\mem_rdata_q[20] ),
    .Y(_14132_));
 sky130_fd_sc_hd__nor3_4 _17753_ (.A(is_alu_reg_imm),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(instr_jalr),
    .Y(_14133_));
 sky130_fd_sc_hd__buf_2 _17754_ (.A(_14133_),
    .X(_14134_));
 sky130_fd_sc_hd__o2bb2ai_1 _17755_ (.A1_N(_14112_),
    .A2_N(\mem_rdata_q[7] ),
    .B1(_14132_),
    .B2(_14134_),
    .Y(_14135_));
 sky130_fd_sc_hd__buf_2 _17756_ (.A(_13005_),
    .X(_14136_));
 sky130_fd_sc_hd__mux2_1 _17757_ (.A0(_14135_),
    .A1(\decoded_imm[0] ),
    .S(_14136_),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_1 _17758_ (.A0(\decoded_rd[4] ),
    .A1(\mem_rdata_latched[11] ),
    .S(_14131_),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_1 _17759_ (.A0(\decoded_rd[3] ),
    .A1(\mem_rdata_latched[10] ),
    .S(_14131_),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_1 _17760_ (.A0(\decoded_rd[2] ),
    .A1(\mem_rdata_latched[9] ),
    .S(_14131_),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_1 _17761_ (.A0(\decoded_rd[1] ),
    .A1(\mem_rdata_latched[8] ),
    .S(_14131_),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_1 _17762_ (.A0(\decoded_rd[0] ),
    .A1(\mem_rdata_latched[7] ),
    .S(_12681_),
    .X(_03179_));
 sky130_fd_sc_hd__buf_1 _17763_ (.A(net494),
    .X(_14137_));
 sky130_fd_sc_hd__buf_2 _17764_ (.A(_14137_),
    .X(_14138_));
 sky130_fd_sc_hd__buf_4 _17765_ (.A(_14138_),
    .X(_14139_));
 sky130_fd_sc_hd__clkbuf_4 _17766_ (.A(_13056_),
    .X(_14140_));
 sky130_fd_sc_hd__buf_4 _17767_ (.A(\mem_rdata_q[27] ),
    .X(_14141_));
 sky130_fd_sc_hd__nand3b_4 _17768_ (.A_N(_13046_),
    .B(_14141_),
    .C(_13048_),
    .Y(_14142_));
 sky130_fd_sc_hd__nand3b_2 _17769_ (.A_N(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[1] ),
    .C(\mem_rdata_q[0] ),
    .Y(_14143_));
 sky130_fd_sc_hd__nor3b_2 _17770_ (.A(\mem_rdata_q[4] ),
    .B(\mem_rdata_q[2] ),
    .C_N(\mem_rdata_q[3] ),
    .Y(_14144_));
 sky130_fd_sc_hd__nor3b_4 _17771_ (.A(\mem_rdata_q[5] ),
    .B(_14143_),
    .C_N(_14144_),
    .Y(_14145_));
 sky130_fd_sc_hd__and3_1 _17772_ (.A(_12996_),
    .B(\mem_rdata_q[25] ),
    .C(_12999_),
    .X(_14146_));
 sky130_fd_sc_hd__nand2_1 _17773_ (.A(_14145_),
    .B(_14146_),
    .Y(_14147_));
 sky130_fd_sc_hd__o2bb2ai_1 _17774_ (.A1_N(_14139_),
    .A2_N(_14140_),
    .B1(_14142_),
    .B2(_14147_),
    .Y(_03178_));
 sky130_fd_sc_hd__nor2_1 _17775_ (.A(_12688_),
    .B(_12690_),
    .Y(_14148_));
 sky130_fd_sc_hd__nand3_1 _17776_ (.A(_14148_),
    .B(\mem_rdata_latched[27] ),
    .C(_12981_),
    .Y(_14149_));
 sky130_fd_sc_hd__o21ai_1 _17777_ (.A1(_12696_),
    .A2(_15210_),
    .B1(_14149_),
    .Y(_03177_));
 sky130_fd_sc_hd__nand3b_1 _17778_ (.A_N(_13046_),
    .B(\mem_rdata_q[26] ),
    .C(_13048_),
    .Y(_14150_));
 sky130_vsdinv _17779_ (.A(\mem_rdata_q[28] ),
    .Y(_14151_));
 sky130_vsdinv _17780_ (.A(_14141_),
    .Y(_14152_));
 sky130_fd_sc_hd__and4b_1 _17781_ (.A_N(_14150_),
    .B(_14145_),
    .C(_14151_),
    .D(_14152_),
    .X(_14153_));
 sky130_fd_sc_hd__buf_2 _17782_ (.A(\mem_rdata_q[25] ),
    .X(_14154_));
 sky130_fd_sc_hd__buf_4 _17783_ (.A(_12955_),
    .X(_14155_));
 sky130_fd_sc_hd__a32o_1 _17784_ (.A1(_14153_),
    .A2(_14154_),
    .A3(_12996_),
    .B1(_14155_),
    .B2(_14122_),
    .X(_03176_));
 sky130_fd_sc_hd__o21ai_1 _17785_ (.A1(_12831_),
    .A2(_15210_),
    .B1(_12695_),
    .Y(_03175_));
 sky130_fd_sc_hd__buf_2 _17786_ (.A(_13059_),
    .X(_14156_));
 sky130_fd_sc_hd__clkbuf_2 _17787_ (.A(_12998_),
    .X(_14157_));
 sky130_fd_sc_hd__and4_1 _17788_ (.A(_14145_),
    .B(_14146_),
    .C(_14152_),
    .D(_14157_),
    .X(_14158_));
 sky130_fd_sc_hd__a21o_1 _17789_ (.A1(instr_setq),
    .A2(_14156_),
    .B1(_14158_),
    .X(_03174_));
 sky130_fd_sc_hd__a22o_1 _17790_ (.A1(instr_getq),
    .A2(_14122_),
    .B1(_13024_),
    .B2(_14145_),
    .X(_03173_));
 sky130_fd_sc_hd__nor3_1 _17791_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .Y(_14159_));
 sky130_fd_sc_hd__or3b_1 _17792_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .C_N(_14159_),
    .X(_14160_));
 sky130_fd_sc_hd__and4_1 _17793_ (.A(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[1] ),
    .D(\mem_rdata_q[0] ),
    .X(_14161_));
 sky130_fd_sc_hd__nor3b_4 _17794_ (.A(\mem_rdata_q[3] ),
    .B(\mem_rdata_q[2] ),
    .C_N(\mem_rdata_q[4] ),
    .Y(_14162_));
 sky130_fd_sc_hd__and3b_1 _17795_ (.A_N(_14160_),
    .B(_14161_),
    .C(_14162_),
    .X(_14163_));
 sky130_vsdinv _17796_ (.A(\mem_rdata_q[23] ),
    .Y(_14164_));
 sky130_vsdinv _17797_ (.A(\mem_rdata_q[22] ),
    .Y(_14165_));
 sky130_fd_sc_hd__nand2_2 _17798_ (.A(_14164_),
    .B(_14165_),
    .Y(_14166_));
 sky130_fd_sc_hd__or4_4 _17799_ (.A(\mem_rdata_q[24] ),
    .B(\mem_rdata_q[21] ),
    .C(\mem_rdata_q[11] ),
    .D(\mem_rdata_q[10] ),
    .X(_14167_));
 sky130_fd_sc_hd__or4b_4 _17800_ (.A(\mem_rdata_q[9] ),
    .B(\mem_rdata_q[8] ),
    .C(\mem_rdata_q[7] ),
    .D_N(_13041_),
    .X(_14168_));
 sky130_fd_sc_hd__nor3_2 _17801_ (.A(_14166_),
    .B(_14167_),
    .C(_14168_),
    .Y(_14169_));
 sky130_fd_sc_hd__a32o_1 _17802_ (.A1(_14163_),
    .A2(_14169_),
    .A3(_13024_),
    .B1(instr_ecall_ebreak),
    .B2(_14122_),
    .X(_03172_));
 sky130_fd_sc_hd__buf_1 _17803_ (.A(instr_rdinstrh),
    .X(_14170_));
 sky130_fd_sc_hd__clkbuf_4 _17804_ (.A(_14170_),
    .X(_14171_));
 sky130_vsdinv _17805_ (.A(\mem_rdata_q[21] ),
    .Y(_14172_));
 sky130_fd_sc_hd__nand3b_4 _17806_ (.A_N(_14166_),
    .B(_14161_),
    .C(_14162_),
    .Y(_14173_));
 sky130_fd_sc_hd__nor3b_4 _17807_ (.A(\mem_rdata_q[20] ),
    .B(_13046_),
    .C_N(_12997_),
    .Y(_14174_));
 sky130_fd_sc_hd__nor3b_4 _17808_ (.A(_14172_),
    .B(_14173_),
    .C_N(_14174_),
    .Y(_14175_));
 sky130_vsdinv _17809_ (.A(_14175_),
    .Y(_14176_));
 sky130_vsdinv _17810_ (.A(\mem_rdata_q[31] ),
    .Y(_14177_));
 sky130_fd_sc_hd__or4_4 _17811_ (.A(\mem_rdata_q[29] ),
    .B(\mem_rdata_q[24] ),
    .C(_14177_),
    .D(_13015_),
    .X(_14178_));
 sky130_fd_sc_hd__or4_4 _17812_ (.A(_13016_),
    .B(_14116_),
    .C(_14178_),
    .D(_14160_),
    .X(_14179_));
 sky130_vsdinv _17813_ (.A(_14154_),
    .Y(_14180_));
 sky130_fd_sc_hd__nand3b_4 _17814_ (.A_N(_14179_),
    .B(_14141_),
    .C(_14180_),
    .Y(_14181_));
 sky130_fd_sc_hd__o2bb2ai_1 _17815_ (.A1_N(_14171_),
    .A2_N(_14140_),
    .B1(_14176_),
    .B2(_14181_),
    .Y(_03171_));
 sky130_fd_sc_hd__buf_2 _17816_ (.A(instr_rdinstr),
    .X(_14182_));
 sky130_fd_sc_hd__buf_4 _17817_ (.A(_14182_),
    .X(_14183_));
 sky130_fd_sc_hd__nand3b_4 _17818_ (.A_N(_14179_),
    .B(_14152_),
    .C(_14180_),
    .Y(_14184_));
 sky130_fd_sc_hd__o2bb2ai_1 _17819_ (.A1_N(_14183_),
    .A2_N(_14140_),
    .B1(_14176_),
    .B2(_14184_),
    .Y(_03170_));
 sky130_fd_sc_hd__buf_2 _17820_ (.A(instr_rdcycleh),
    .X(_14185_));
 sky130_fd_sc_hd__clkbuf_4 _17821_ (.A(_14185_),
    .X(_14186_));
 sky130_fd_sc_hd__nor3_4 _17822_ (.A(\mem_rdata_q[21] ),
    .B(_13005_),
    .C(_14173_),
    .Y(_14187_));
 sky130_vsdinv _17823_ (.A(_14187_),
    .Y(_14188_));
 sky130_fd_sc_hd__o2bb2ai_1 _17824_ (.A1_N(_14186_),
    .A2_N(_14140_),
    .B1(_14188_),
    .B2(_14181_),
    .Y(_03169_));
 sky130_fd_sc_hd__o2bb2ai_1 _17825_ (.A1_N(instr_rdcycle),
    .A2_N(_14140_),
    .B1(_14188_),
    .B2(_14184_),
    .Y(_03168_));
 sky130_fd_sc_hd__nor3b_4 _17826_ (.A(_13014_),
    .B(_13046_),
    .C_N(_13048_),
    .Y(_14189_));
 sky130_fd_sc_hd__nand3b_1 _17827_ (.A_N(_13017_),
    .B(_13021_),
    .C(_14189_),
    .Y(_14190_));
 sky130_fd_sc_hd__o2bb2ai_1 _17828_ (.A1_N(instr_srai),
    .A2_N(_14140_),
    .B1(_14102_),
    .B2(_14190_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand3_1 _17829_ (.A(_13024_),
    .B(_13047_),
    .C(_13021_),
    .Y(_14191_));
 sky130_fd_sc_hd__o21ai_1 _17830_ (.A1(_12827_),
    .A2(_14113_),
    .B1(_14191_),
    .Y(_03166_));
 sky130_fd_sc_hd__a32o_1 _17831_ (.A1(_13024_),
    .A2(_13047_),
    .A3(_13038_),
    .B1(instr_slli),
    .B2(_14122_),
    .X(_03165_));
 sky130_fd_sc_hd__and2_1 _17832_ (.A(_13033_),
    .B(_14157_),
    .X(_14192_));
 sky130_fd_sc_hd__a22o_1 _17833_ (.A1(instr_sw),
    .A2(_14122_),
    .B1(_14192_),
    .B2(_14112_),
    .X(_03164_));
 sky130_fd_sc_hd__and2_1 _17834_ (.A(_13038_),
    .B(_14157_),
    .X(_14193_));
 sky130_fd_sc_hd__a22o_1 _17835_ (.A1(instr_sh),
    .A2(_13060_),
    .B1(_14193_),
    .B2(_14112_),
    .X(_03163_));
 sky130_fd_sc_hd__and2_1 _17836_ (.A(_13041_),
    .B(_14157_),
    .X(_14194_));
 sky130_fd_sc_hd__a22o_1 _17837_ (.A1(instr_sb),
    .A2(_13060_),
    .B1(_14194_),
    .B2(_14112_),
    .X(_03162_));
 sky130_vsdinv _17838_ (.A(instr_lhu),
    .Y(_14195_));
 sky130_fd_sc_hd__buf_2 _17839_ (.A(_14157_),
    .X(_14196_));
 sky130_fd_sc_hd__nand3b_1 _17840_ (.A_N(_13020_),
    .B(_14123_),
    .C(_14196_),
    .Y(_14197_));
 sky130_fd_sc_hd__o21ai_1 _17841_ (.A1(_14195_),
    .A2(_14113_),
    .B1(_14197_),
    .Y(_03161_));
 sky130_fd_sc_hd__nand3_1 _17842_ (.A(_13027_),
    .B(_14123_),
    .C(_14196_),
    .Y(_14198_));
 sky130_fd_sc_hd__a21bo_1 _17843_ (.A1(instr_lbu),
    .A2(_14156_),
    .B1_N(_14198_),
    .X(_03160_));
 sky130_fd_sc_hd__a22o_1 _17844_ (.A1(instr_lw),
    .A2(_13060_),
    .B1(_14192_),
    .B2(_14123_),
    .X(_03159_));
 sky130_fd_sc_hd__o2bb2ai_1 _17845_ (.A1_N(_14123_),
    .A2_N(_14193_),
    .B1(_12657_),
    .B2(_14113_),
    .Y(_03158_));
 sky130_fd_sc_hd__a22o_1 _17846_ (.A1(instr_lb),
    .A2(_13060_),
    .B1(_14194_),
    .B2(_14123_),
    .X(_03157_));
 sky130_fd_sc_hd__nand3_2 _17847_ (.A(_00325_),
    .B(_00324_),
    .C(_00326_),
    .Y(_14199_));
 sky130_fd_sc_hd__or2b_1 _17848_ (.A(_14199_),
    .B_N(_12682_),
    .X(_14200_));
 sky130_fd_sc_hd__or4_4 _17849_ (.A(\mem_rdata_latched[14] ),
    .B(\mem_rdata_latched[13] ),
    .C(\mem_rdata_latched[12] ),
    .D(_12982_),
    .X(_14201_));
 sky130_fd_sc_hd__nor3b_2 _17850_ (.A(_14200_),
    .B(_14201_),
    .C_N(_12681_),
    .Y(_14202_));
 sky130_fd_sc_hd__a21o_1 _17851_ (.A1(instr_jalr),
    .A2(_00337_),
    .B1(_14202_),
    .X(_03156_));
 sky130_fd_sc_hd__or4_4 _17852_ (.A(_12682_),
    .B(_12982_),
    .C(_14199_),
    .D(_12692_),
    .X(_14203_));
 sky130_fd_sc_hd__o21ai_1 _17853_ (.A1(_00323_),
    .A2(_15210_),
    .B1(_14203_),
    .Y(_03155_));
 sky130_fd_sc_hd__and4b_1 _17854_ (.A_N(_14200_),
    .B(_14100_),
    .C(_00328_),
    .D(_12686_),
    .X(_14204_));
 sky130_fd_sc_hd__a22o_1 _17855_ (.A1(instr_auipc),
    .A2(_12984_),
    .B1(_14204_),
    .B2(_12684_),
    .X(_03154_));
 sky130_fd_sc_hd__clkbuf_4 _17856_ (.A(instr_lui),
    .X(_14205_));
 sky130_fd_sc_hd__a22o_1 _17857_ (.A1(_14205_),
    .A2(_12984_),
    .B1(_14204_),
    .B2(_00329_),
    .X(_03153_));
 sky130_fd_sc_hd__clkbuf_2 _17858_ (.A(\mem_rdata_q[31] ),
    .X(_14206_));
 sky130_fd_sc_hd__buf_2 _17859_ (.A(_14206_),
    .X(_14207_));
 sky130_fd_sc_hd__mux2_1 _17860_ (.A0(net298),
    .A1(_14207_),
    .S(_14196_),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_1 _17861_ (.A0(net297),
    .A1(\mem_rdata_q[30] ),
    .S(_14196_),
    .X(_03151_));
 sky130_fd_sc_hd__o21ba_1 _17862_ (.A1(net295),
    .A2(_13572_),
    .B1_N(_14189_),
    .X(_03150_));
 sky130_fd_sc_hd__mux2_1 _17863_ (.A0(net294),
    .A1(\mem_rdata_q[28] ),
    .S(_14196_),
    .X(_03149_));
 sky130_fd_sc_hd__a21bo_1 _17864_ (.A1(_14156_),
    .A2(net293),
    .B1_N(_14142_),
    .X(_03148_));
 sky130_fd_sc_hd__a21bo_1 _17865_ (.A1(_14156_),
    .A2(net292),
    .B1_N(_14150_),
    .X(_03147_));
 sky130_fd_sc_hd__mux2_1 _17866_ (.A0(net291),
    .A1(_14154_),
    .S(_14196_),
    .X(_03146_));
 sky130_fd_sc_hd__buf_2 _17867_ (.A(_13062_),
    .X(_14208_));
 sky130_fd_sc_hd__mux2_1 _17868_ (.A0(net290),
    .A1(\mem_rdata_q[24] ),
    .S(_14208_),
    .X(_03145_));
 sky130_fd_sc_hd__mux2_1 _17869_ (.A0(net289),
    .A1(\mem_rdata_q[23] ),
    .S(_14208_),
    .X(_03144_));
 sky130_fd_sc_hd__mux2_1 _17870_ (.A0(net288),
    .A1(\mem_rdata_q[22] ),
    .S(_14208_),
    .X(_03143_));
 sky130_fd_sc_hd__mux2_1 _17871_ (.A0(net287),
    .A1(\mem_rdata_q[21] ),
    .S(_14208_),
    .X(_03142_));
 sky130_fd_sc_hd__o21ba_1 _17872_ (.A1(net286),
    .A2(_13572_),
    .B1_N(_14174_),
    .X(_03141_));
 sky130_fd_sc_hd__mux2_1 _17873_ (.A0(net284),
    .A1(\mem_rdata_q[19] ),
    .S(_14208_),
    .X(_03140_));
 sky130_fd_sc_hd__mux2_1 _17874_ (.A0(net283),
    .A1(\mem_rdata_q[18] ),
    .S(_14208_),
    .X(_03139_));
 sky130_fd_sc_hd__clkbuf_4 _17875_ (.A(_13062_),
    .X(_14209_));
 sky130_fd_sc_hd__mux2_1 _17876_ (.A0(net282),
    .A1(\mem_rdata_q[17] ),
    .S(_14209_),
    .X(_03138_));
 sky130_fd_sc_hd__mux2_1 _17877_ (.A0(net281),
    .A1(\mem_rdata_q[16] ),
    .S(_14209_),
    .X(_03137_));
 sky130_fd_sc_hd__mux2_1 _17878_ (.A0(net280),
    .A1(\mem_rdata_q[15] ),
    .S(_14209_),
    .X(_03136_));
 sky130_fd_sc_hd__mux2_1 _17879_ (.A0(net279),
    .A1(_12990_),
    .S(_14209_),
    .X(_03135_));
 sky130_fd_sc_hd__mux2_1 _17880_ (.A0(net278),
    .A1(_12992_),
    .S(_14209_),
    .X(_03134_));
 sky130_fd_sc_hd__mux2_1 _17881_ (.A0(net277),
    .A1(_12994_),
    .S(_14209_),
    .X(_03133_));
 sky130_fd_sc_hd__buf_2 _17882_ (.A(_13062_),
    .X(_14210_));
 sky130_fd_sc_hd__mux2_1 _17883_ (.A0(net276),
    .A1(\mem_rdata_q[11] ),
    .S(_14210_),
    .X(_03132_));
 sky130_fd_sc_hd__mux2_1 _17884_ (.A0(net275),
    .A1(\mem_rdata_q[10] ),
    .S(_14210_),
    .X(_03131_));
 sky130_fd_sc_hd__mux2_1 _17885_ (.A0(net305),
    .A1(\mem_rdata_q[9] ),
    .S(_14210_),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_1 _17886_ (.A0(net304),
    .A1(\mem_rdata_q[8] ),
    .S(_14210_),
    .X(_03129_));
 sky130_fd_sc_hd__mux2_1 _17887_ (.A0(net303),
    .A1(\mem_rdata_q[7] ),
    .S(_14210_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_1 _17888_ (.A0(net302),
    .A1(\mem_rdata_q[6] ),
    .S(_14210_),
    .X(_03127_));
 sky130_fd_sc_hd__buf_2 _17889_ (.A(_13062_),
    .X(_14211_));
 sky130_fd_sc_hd__mux2_1 _17890_ (.A0(net301),
    .A1(\mem_rdata_q[5] ),
    .S(_14211_),
    .X(_03126_));
 sky130_fd_sc_hd__mux2_1 _17891_ (.A0(net300),
    .A1(\mem_rdata_q[4] ),
    .S(_14211_),
    .X(_03125_));
 sky130_fd_sc_hd__mux2_1 _17892_ (.A0(net299),
    .A1(\mem_rdata_q[3] ),
    .S(_14211_),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_1 _17893_ (.A0(net296),
    .A1(\mem_rdata_q[2] ),
    .S(_14211_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_1 _17894_ (.A0(net285),
    .A1(\mem_rdata_q[1] ),
    .S(_14211_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_1 _17895_ (.A0(net274),
    .A1(\mem_rdata_q[0] ),
    .S(_14211_),
    .X(_03121_));
 sky130_fd_sc_hd__buf_2 _17896_ (.A(\cpu_state[5] ),
    .X(_14212_));
 sky130_fd_sc_hd__nor3_1 _17897_ (.A(_12849_),
    .B(_12651_),
    .C(_14212_),
    .Y(_14213_));
 sky130_fd_sc_hd__or4_4 _17898_ (.A(_12642_),
    .B(_00318_),
    .C(_00320_),
    .D(_14213_),
    .X(_14214_));
 sky130_fd_sc_hd__buf_4 _17899_ (.A(_14214_),
    .X(_14215_));
 sky130_fd_sc_hd__buf_2 _17900_ (.A(_14215_),
    .X(_14216_));
 sky130_fd_sc_hd__mux2_1 _17901_ (.A0(_02499_),
    .A1(_12797_),
    .S(_14216_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_4 _17902_ (.A(net329),
    .X(_14217_));
 sky130_fd_sc_hd__mux2_1 _17903_ (.A0(_02498_),
    .A1(_14217_),
    .S(_14216_),
    .X(_03119_));
 sky130_fd_sc_hd__buf_2 _17904_ (.A(net327),
    .X(_14218_));
 sky130_fd_sc_hd__mux2_1 _17905_ (.A0(_02496_),
    .A1(_14218_),
    .S(_14216_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_2 _17906_ (.A(net326),
    .X(_14219_));
 sky130_fd_sc_hd__clkbuf_4 _17907_ (.A(_14219_),
    .X(_14220_));
 sky130_fd_sc_hd__mux2_1 _17908_ (.A0(_02495_),
    .A1(_14220_),
    .S(_14216_),
    .X(_03117_));
 sky130_fd_sc_hd__clkbuf_2 _17909_ (.A(net325),
    .X(_14221_));
 sky130_fd_sc_hd__buf_2 _17910_ (.A(_14221_),
    .X(_14222_));
 sky130_fd_sc_hd__mux2_1 _17911_ (.A0(_02494_),
    .A1(_14222_),
    .S(_14216_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_4 _17912_ (.A(net324),
    .X(_14223_));
 sky130_fd_sc_hd__buf_2 _17913_ (.A(_14223_),
    .X(_14224_));
 sky130_fd_sc_hd__mux2_1 _17914_ (.A0(_02493_),
    .A1(_14224_),
    .S(_14216_),
    .X(_03115_));
 sky130_fd_sc_hd__buf_2 _17915_ (.A(net323),
    .X(_14225_));
 sky130_fd_sc_hd__clkbuf_4 _17916_ (.A(_14225_),
    .X(_14226_));
 sky130_fd_sc_hd__buf_2 _17917_ (.A(_14215_),
    .X(_14227_));
 sky130_fd_sc_hd__mux2_1 _17918_ (.A0(_02492_),
    .A1(_14226_),
    .S(_14227_),
    .X(_03114_));
 sky130_fd_sc_hd__buf_4 _17919_ (.A(net322),
    .X(_14228_));
 sky130_fd_sc_hd__clkbuf_4 _17920_ (.A(_14228_),
    .X(_14229_));
 sky130_fd_sc_hd__mux2_1 _17921_ (.A0(_02491_),
    .A1(_14229_),
    .S(_14227_),
    .X(_03113_));
 sky130_fd_sc_hd__clkbuf_4 _17922_ (.A(net321),
    .X(_14230_));
 sky130_fd_sc_hd__mux2_1 _17923_ (.A0(_02490_),
    .A1(_14230_),
    .S(_14227_),
    .X(_03112_));
 sky130_fd_sc_hd__buf_4 _17924_ (.A(net320),
    .X(_14231_));
 sky130_fd_sc_hd__mux2_1 _17925_ (.A0(_02489_),
    .A1(_14231_),
    .S(_14227_),
    .X(_03111_));
 sky130_fd_sc_hd__buf_4 _17926_ (.A(net319),
    .X(_14232_));
 sky130_fd_sc_hd__mux2_1 _17927_ (.A0(_02488_),
    .A1(_14232_),
    .S(_14227_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_4 _17928_ (.A(net318),
    .X(_14233_));
 sky130_fd_sc_hd__mux2_1 _17929_ (.A0(_02487_),
    .A1(_14233_),
    .S(_14227_),
    .X(_03109_));
 sky130_fd_sc_hd__buf_4 _17930_ (.A(net316),
    .X(_14234_));
 sky130_fd_sc_hd__buf_2 _17931_ (.A(_14215_),
    .X(_14235_));
 sky130_fd_sc_hd__mux2_1 _17932_ (.A0(_02485_),
    .A1(_14234_),
    .S(_14235_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_4 _17933_ (.A(net315),
    .X(_14236_));
 sky130_fd_sc_hd__mux2_1 _17934_ (.A0(_02484_),
    .A1(_14236_),
    .S(_14235_),
    .X(_03107_));
 sky130_fd_sc_hd__buf_2 _17935_ (.A(net314),
    .X(_14237_));
 sky130_fd_sc_hd__buf_4 _17936_ (.A(_14237_),
    .X(_14238_));
 sky130_fd_sc_hd__mux2_1 _17937_ (.A0(_02483_),
    .A1(_14238_),
    .S(_14235_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_4 _17938_ (.A(net313),
    .X(_14239_));
 sky130_fd_sc_hd__buf_4 _17939_ (.A(_14239_),
    .X(_14240_));
 sky130_fd_sc_hd__mux2_1 _17940_ (.A0(_02482_),
    .A1(_14240_),
    .S(_14235_),
    .X(_03105_));
 sky130_fd_sc_hd__buf_6 _17941_ (.A(net312),
    .X(_14241_));
 sky130_fd_sc_hd__mux2_1 _17942_ (.A0(_02481_),
    .A1(_14241_),
    .S(_14235_),
    .X(_03104_));
 sky130_fd_sc_hd__buf_6 _17943_ (.A(net311),
    .X(_14242_));
 sky130_fd_sc_hd__mux2_1 _17944_ (.A0(_02480_),
    .A1(_14242_),
    .S(_14235_),
    .X(_03103_));
 sky130_fd_sc_hd__buf_6 _17945_ (.A(net310),
    .X(_14243_));
 sky130_fd_sc_hd__buf_2 _17946_ (.A(_14215_),
    .X(_14244_));
 sky130_fd_sc_hd__mux2_1 _17947_ (.A0(_02479_),
    .A1(_14243_),
    .S(_14244_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_6 _17948_ (.A(net309),
    .X(_14245_));
 sky130_fd_sc_hd__mux2_1 _17949_ (.A0(_02478_),
    .A1(_14245_),
    .S(_14244_),
    .X(_03101_));
 sky130_fd_sc_hd__clkbuf_8 _17950_ (.A(net308),
    .X(_14246_));
 sky130_fd_sc_hd__mux2_1 _17951_ (.A0(_02477_),
    .A1(_14246_),
    .S(_14244_),
    .X(_03100_));
 sky130_fd_sc_hd__buf_6 _17952_ (.A(net307),
    .X(_14247_));
 sky130_fd_sc_hd__mux2_1 _17953_ (.A0(_02476_),
    .A1(_14247_),
    .S(_14244_),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_4 _17954_ (.A(net337),
    .X(_14248_));
 sky130_fd_sc_hd__buf_4 _17955_ (.A(_14248_),
    .X(_14249_));
 sky130_fd_sc_hd__mux2_1 _17956_ (.A0(_02506_),
    .A1(_14249_),
    .S(_14244_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_4 _17957_ (.A(net336),
    .X(_14250_));
 sky130_fd_sc_hd__buf_6 _17958_ (.A(_14250_),
    .X(_14251_));
 sky130_fd_sc_hd__mux2_1 _17959_ (.A0(_02505_),
    .A1(_14251_),
    .S(_14244_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_4 _17960_ (.A(net335),
    .X(_14252_));
 sky130_fd_sc_hd__buf_4 _17961_ (.A(_14252_),
    .X(_14253_));
 sky130_fd_sc_hd__clkbuf_4 _17962_ (.A(_14214_),
    .X(_14254_));
 sky130_fd_sc_hd__mux2_1 _17963_ (.A0(_02504_),
    .A1(_14253_),
    .S(_14254_),
    .X(_03096_));
 sky130_fd_sc_hd__buf_4 _17964_ (.A(net334),
    .X(_14255_));
 sky130_fd_sc_hd__buf_4 _17965_ (.A(_14255_),
    .X(_14256_));
 sky130_fd_sc_hd__mux2_1 _17966_ (.A0(_02503_),
    .A1(_14256_),
    .S(_14254_),
    .X(_03095_));
 sky130_fd_sc_hd__buf_6 _17967_ (.A(net333),
    .X(_14257_));
 sky130_fd_sc_hd__mux2_1 _17968_ (.A0(_02502_),
    .A1(_14257_),
    .S(_14254_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_4 _17969_ (.A(net332),
    .X(_14258_));
 sky130_fd_sc_hd__buf_6 _17970_ (.A(_14258_),
    .X(_14259_));
 sky130_fd_sc_hd__mux2_1 _17971_ (.A0(_02501_),
    .A1(_14259_),
    .S(_14254_),
    .X(_03093_));
 sky130_fd_sc_hd__buf_4 _17972_ (.A(net331),
    .X(_14260_));
 sky130_fd_sc_hd__mux2_1 _17973_ (.A0(_02500_),
    .A1(_14260_),
    .S(_14254_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_4 _17974_ (.A(net328),
    .X(_14261_));
 sky130_fd_sc_hd__buf_6 _17975_ (.A(_14261_),
    .X(_14262_));
 sky130_fd_sc_hd__mux2_1 _17976_ (.A0(_02497_),
    .A1(_14262_),
    .S(_14254_),
    .X(_03091_));
 sky130_fd_sc_hd__buf_6 _17977_ (.A(net317),
    .X(_14263_));
 sky130_fd_sc_hd__clkbuf_2 _17978_ (.A(_14263_),
    .X(_14264_));
 sky130_fd_sc_hd__buf_2 _17979_ (.A(_14264_),
    .X(_14265_));
 sky130_fd_sc_hd__mux2_1 _17980_ (.A0(_02486_),
    .A1(_14265_),
    .S(_14215_),
    .X(_03090_));
 sky130_fd_sc_hd__buf_4 _17981_ (.A(net306),
    .X(_14266_));
 sky130_fd_sc_hd__buf_6 _17982_ (.A(_14266_),
    .X(_14267_));
 sky130_fd_sc_hd__clkbuf_2 _17983_ (.A(_14267_),
    .X(_14268_));
 sky130_fd_sc_hd__buf_2 _17984_ (.A(_14268_),
    .X(_14269_));
 sky130_fd_sc_hd__mux2_1 _17985_ (.A0(_02475_),
    .A1(_14269_),
    .S(_14215_),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_1 _17986_ (.A0(net191),
    .A1(net158),
    .S(net431),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_1 _17987_ (.A0(net190),
    .A1(net157),
    .S(_12975_),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_1 _17988_ (.A0(net188),
    .A1(net155),
    .S(net431),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_1 _17989_ (.A0(net187),
    .A1(net154),
    .S(net431),
    .X(_03085_));
 sky130_fd_sc_hd__mux2_1 _17990_ (.A0(net186),
    .A1(net153),
    .S(_12975_),
    .X(_03084_));
 sky130_fd_sc_hd__clkbuf_4 _17991_ (.A(_12974_),
    .X(_14270_));
 sky130_fd_sc_hd__mux2_1 _17992_ (.A0(net185),
    .A1(net152),
    .S(net430),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_1 _17993_ (.A0(net184),
    .A1(net151),
    .S(net430),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_1 _17994_ (.A0(net183),
    .A1(net150),
    .S(net430),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_1 _17995_ (.A0(net182),
    .A1(net149),
    .S(net430),
    .X(_03080_));
 sky130_fd_sc_hd__mux2_1 _17996_ (.A0(net181),
    .A1(net148),
    .S(_14270_),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_1 _17997_ (.A0(net180),
    .A1(net147),
    .S(net430),
    .X(_03078_));
 sky130_fd_sc_hd__buf_6 _17998_ (.A(_12974_),
    .X(_14271_));
 sky130_fd_sc_hd__mux2_1 _17999_ (.A0(net179),
    .A1(net146),
    .S(net429),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_1 _18000_ (.A0(net177),
    .A1(net144),
    .S(net429),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_1 _18001_ (.A0(net176),
    .A1(net143),
    .S(net429),
    .X(_03075_));
 sky130_fd_sc_hd__mux2_1 _18002_ (.A0(net175),
    .A1(net142),
    .S(_14271_),
    .X(_03074_));
 sky130_fd_sc_hd__mux2_1 _18003_ (.A0(net174),
    .A1(net141),
    .S(_14271_),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_1 _18004_ (.A0(net173),
    .A1(net140),
    .S(net429),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_2 _18005_ (.A(_12974_),
    .X(_14272_));
 sky130_fd_sc_hd__mux2_1 _18006_ (.A0(net172),
    .A1(net139),
    .S(net428),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_1 _18007_ (.A0(net171),
    .A1(net138),
    .S(net427),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _18008_ (.A0(net170),
    .A1(net137),
    .S(net427),
    .X(_03069_));
 sky130_fd_sc_hd__mux2_1 _18009_ (.A0(net169),
    .A1(net136),
    .S(net427),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_1 _18010_ (.A0(net168),
    .A1(net135),
    .S(_14272_),
    .X(_03067_));
 sky130_fd_sc_hd__mux2_1 _18011_ (.A0(net198),
    .A1(net165),
    .S(net428),
    .X(_03066_));
 sky130_fd_sc_hd__buf_6 _18012_ (.A(_12974_),
    .X(_14273_));
 sky130_fd_sc_hd__mux2_1 _18013_ (.A0(net197),
    .A1(net164),
    .S(_14273_),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_1 _18014_ (.A0(net196),
    .A1(net163),
    .S(_14273_),
    .X(_03064_));
 sky130_fd_sc_hd__mux2_1 _18015_ (.A0(net195),
    .A1(net162),
    .S(_14273_),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_1 _18016_ (.A0(net194),
    .A1(net161),
    .S(_14273_),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_1 _18017_ (.A0(net193),
    .A1(net160),
    .S(_14273_),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_1 _18018_ (.A0(net192),
    .A1(net159),
    .S(_14273_),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_1 _18019_ (.A0(net189),
    .A1(net156),
    .S(_12974_),
    .X(_03059_));
 sky130_vsdinv _18020_ (.A(\pcpi_mul.rs1[31] ),
    .Y(_14274_));
 sky130_fd_sc_hd__buf_4 _18021_ (.A(_14274_),
    .X(_14275_));
 sky130_fd_sc_hd__buf_6 _18022_ (.A(_14275_),
    .X(_14276_));
 sky130_fd_sc_hd__buf_6 _18023_ (.A(_14276_),
    .X(_14277_));
 sky130_fd_sc_hd__o21ai_1 _18024_ (.A1(_14277_),
    .A2(_14079_),
    .B1(_12798_),
    .Y(_03058_));
 sky130_vsdinv _18025_ (.A(\pcpi_mul.rs1[30] ),
    .Y(_14278_));
 sky130_fd_sc_hd__clkbuf_4 _18026_ (.A(_14278_),
    .X(_14279_));
 sky130_fd_sc_hd__buf_4 _18027_ (.A(_14279_),
    .X(_14280_));
 sky130_fd_sc_hd__buf_6 _18028_ (.A(_14280_),
    .X(_14281_));
 sky130_fd_sc_hd__clkbuf_2 _18029_ (.A(_14078_),
    .X(_14282_));
 sky130_fd_sc_hd__nand2_1 _18030_ (.A(_14080_),
    .B(_14217_),
    .Y(_14283_));
 sky130_fd_sc_hd__o21ai_1 _18031_ (.A1(_14281_),
    .A2(_14282_),
    .B1(_14283_),
    .Y(_03057_));
 sky130_vsdinv _18032_ (.A(\pcpi_mul.rs1[29] ),
    .Y(_14284_));
 sky130_fd_sc_hd__buf_2 _18033_ (.A(_14284_),
    .X(_14285_));
 sky130_fd_sc_hd__buf_4 _18034_ (.A(_14285_),
    .X(_14286_));
 sky130_fd_sc_hd__buf_6 _18035_ (.A(_14286_),
    .X(_14287_));
 sky130_fd_sc_hd__clkbuf_2 _18036_ (.A(_12793_),
    .X(_14288_));
 sky130_fd_sc_hd__nand2_1 _18037_ (.A(_14288_),
    .B(_14218_),
    .Y(_14289_));
 sky130_fd_sc_hd__o21ai_1 _18038_ (.A1(_14287_),
    .A2(_14282_),
    .B1(_14289_),
    .Y(_03056_));
 sky130_vsdinv _18039_ (.A(\pcpi_mul.rs1[28] ),
    .Y(_14290_));
 sky130_fd_sc_hd__buf_4 _18040_ (.A(_14290_),
    .X(_14291_));
 sky130_fd_sc_hd__buf_6 _18041_ (.A(_14291_),
    .X(_14292_));
 sky130_fd_sc_hd__clkbuf_8 _18042_ (.A(_14292_),
    .X(_14293_));
 sky130_fd_sc_hd__buf_6 _18043_ (.A(_14293_),
    .X(_14294_));
 sky130_fd_sc_hd__nand2_1 _18044_ (.A(_14288_),
    .B(_14220_),
    .Y(_14295_));
 sky130_fd_sc_hd__o21ai_1 _18045_ (.A1(_14294_),
    .A2(_14282_),
    .B1(_14295_),
    .Y(_03055_));
 sky130_vsdinv _18046_ (.A(\pcpi_mul.rs1[27] ),
    .Y(_14296_));
 sky130_fd_sc_hd__buf_4 _18047_ (.A(_14296_),
    .X(_14297_));
 sky130_fd_sc_hd__buf_6 _18048_ (.A(_14297_),
    .X(_14298_));
 sky130_fd_sc_hd__clkbuf_8 _18049_ (.A(_14298_),
    .X(_14299_));
 sky130_fd_sc_hd__buf_6 _18050_ (.A(_14299_),
    .X(_14300_));
 sky130_fd_sc_hd__nand2_1 _18051_ (.A(_14288_),
    .B(_14222_),
    .Y(_14301_));
 sky130_fd_sc_hd__o21ai_1 _18052_ (.A1(_14300_),
    .A2(_14282_),
    .B1(_14301_),
    .Y(_03054_));
 sky130_vsdinv _18053_ (.A(\pcpi_mul.rs1[26] ),
    .Y(_14302_));
 sky130_fd_sc_hd__buf_4 _18054_ (.A(_14302_),
    .X(_14303_));
 sky130_fd_sc_hd__buf_4 _18055_ (.A(_14303_),
    .X(_14304_));
 sky130_fd_sc_hd__buf_6 _18056_ (.A(_14304_),
    .X(_14305_));
 sky130_fd_sc_hd__nand2_1 _18057_ (.A(_14288_),
    .B(_14224_),
    .Y(_14306_));
 sky130_fd_sc_hd__o21ai_1 _18058_ (.A1(_14305_),
    .A2(_14282_),
    .B1(_14306_),
    .Y(_03053_));
 sky130_vsdinv _18059_ (.A(\pcpi_mul.rs1[25] ),
    .Y(_14307_));
 sky130_fd_sc_hd__clkbuf_4 _18060_ (.A(_14307_),
    .X(_14308_));
 sky130_fd_sc_hd__buf_4 _18061_ (.A(_14308_),
    .X(_14309_));
 sky130_fd_sc_hd__buf_6 _18062_ (.A(_14309_),
    .X(_14310_));
 sky130_fd_sc_hd__buf_6 _18063_ (.A(_14310_),
    .X(_14311_));
 sky130_fd_sc_hd__nand2_1 _18064_ (.A(_14288_),
    .B(_14226_),
    .Y(_14312_));
 sky130_fd_sc_hd__o21ai_1 _18065_ (.A1(_14311_),
    .A2(_14282_),
    .B1(_14312_),
    .Y(_03052_));
 sky130_vsdinv _18066_ (.A(\pcpi_mul.rs1[24] ),
    .Y(_14313_));
 sky130_fd_sc_hd__buf_4 _18067_ (.A(_14313_),
    .X(_14314_));
 sky130_fd_sc_hd__buf_4 _18068_ (.A(_14314_),
    .X(_14315_));
 sky130_fd_sc_hd__buf_6 _18069_ (.A(_14315_),
    .X(_14316_));
 sky130_fd_sc_hd__clkbuf_2 _18070_ (.A(_14078_),
    .X(_14317_));
 sky130_fd_sc_hd__nand2_1 _18071_ (.A(_14288_),
    .B(_14229_),
    .Y(_14318_));
 sky130_fd_sc_hd__o21ai_1 _18072_ (.A1(_14316_),
    .A2(_14317_),
    .B1(_14318_),
    .Y(_03051_));
 sky130_vsdinv _18073_ (.A(\pcpi_mul.rs1[23] ),
    .Y(_14319_));
 sky130_fd_sc_hd__buf_4 _18074_ (.A(_14319_),
    .X(_14320_));
 sky130_fd_sc_hd__buf_6 _18075_ (.A(_14320_),
    .X(_14321_));
 sky130_fd_sc_hd__buf_6 _18076_ (.A(_14321_),
    .X(_14322_));
 sky130_fd_sc_hd__clkbuf_2 _18077_ (.A(_12795_),
    .X(_14323_));
 sky130_fd_sc_hd__nand2_1 _18078_ (.A(_14323_),
    .B(_14230_),
    .Y(_14324_));
 sky130_fd_sc_hd__o21ai_1 _18079_ (.A1(_14322_),
    .A2(_14317_),
    .B1(_14324_),
    .Y(_03050_));
 sky130_fd_sc_hd__buf_2 _18080_ (.A(\pcpi_mul.rs1[22] ),
    .X(_14325_));
 sky130_vsdinv _18081_ (.A(_14325_),
    .Y(_14326_));
 sky130_fd_sc_hd__buf_4 _18082_ (.A(_14326_),
    .X(_14327_));
 sky130_fd_sc_hd__buf_6 _18083_ (.A(_14327_),
    .X(_14328_));
 sky130_fd_sc_hd__buf_6 _18084_ (.A(_14328_),
    .X(_14329_));
 sky130_fd_sc_hd__nand2_1 _18085_ (.A(_14323_),
    .B(_14231_),
    .Y(_14330_));
 sky130_fd_sc_hd__o21ai_1 _18086_ (.A1(_14329_),
    .A2(_14317_),
    .B1(_14330_),
    .Y(_03049_));
 sky130_fd_sc_hd__clkbuf_4 _18087_ (.A(\pcpi_mul.rs1[21] ),
    .X(_14331_));
 sky130_vsdinv _18088_ (.A(_14331_),
    .Y(_14332_));
 sky130_fd_sc_hd__buf_6 _18089_ (.A(_14332_),
    .X(_14333_));
 sky130_fd_sc_hd__clkbuf_8 _18090_ (.A(_14333_),
    .X(_14334_));
 sky130_fd_sc_hd__buf_6 _18091_ (.A(_14334_),
    .X(_14335_));
 sky130_fd_sc_hd__nand2_1 _18092_ (.A(_14323_),
    .B(_14232_),
    .Y(_14336_));
 sky130_fd_sc_hd__o21ai_1 _18093_ (.A1(_14335_),
    .A2(_14317_),
    .B1(_14336_),
    .Y(_03048_));
 sky130_fd_sc_hd__buf_2 _18094_ (.A(\pcpi_mul.rs1[20] ),
    .X(_14337_));
 sky130_vsdinv _18095_ (.A(_14337_),
    .Y(_14338_));
 sky130_fd_sc_hd__buf_6 _18096_ (.A(_14338_),
    .X(_14339_));
 sky130_fd_sc_hd__buf_6 _18097_ (.A(_14339_),
    .X(_14340_));
 sky130_fd_sc_hd__buf_6 _18098_ (.A(_14340_),
    .X(_14341_));
 sky130_fd_sc_hd__clkbuf_8 _18099_ (.A(_14341_),
    .X(_14342_));
 sky130_fd_sc_hd__nand2_1 _18100_ (.A(_14323_),
    .B(_14233_),
    .Y(_14343_));
 sky130_fd_sc_hd__o21ai_1 _18101_ (.A1(_14342_),
    .A2(_14317_),
    .B1(_14343_),
    .Y(_03047_));
 sky130_fd_sc_hd__clkbuf_4 _18102_ (.A(\pcpi_mul.rs1[19] ),
    .X(_14344_));
 sky130_vsdinv _18103_ (.A(_14344_),
    .Y(_14345_));
 sky130_fd_sc_hd__clkbuf_4 _18104_ (.A(_14345_),
    .X(_14346_));
 sky130_fd_sc_hd__buf_6 _18105_ (.A(_14346_),
    .X(_14347_));
 sky130_fd_sc_hd__buf_6 _18106_ (.A(_14347_),
    .X(_14348_));
 sky130_fd_sc_hd__nand2_1 _18107_ (.A(_14323_),
    .B(_14234_),
    .Y(_14349_));
 sky130_fd_sc_hd__o21ai_1 _18108_ (.A1(_14348_),
    .A2(_14317_),
    .B1(_14349_),
    .Y(_03046_));
 sky130_fd_sc_hd__buf_2 _18109_ (.A(\pcpi_mul.rs1[18] ),
    .X(_14350_));
 sky130_vsdinv _18110_ (.A(_14350_),
    .Y(_14351_));
 sky130_fd_sc_hd__buf_4 _18111_ (.A(_14351_),
    .X(_14352_));
 sky130_fd_sc_hd__buf_4 _18112_ (.A(_14352_),
    .X(_14353_));
 sky130_fd_sc_hd__buf_6 _18113_ (.A(_14353_),
    .X(_14354_));
 sky130_fd_sc_hd__clkbuf_2 _18114_ (.A(_14078_),
    .X(_14355_));
 sky130_fd_sc_hd__nand2_1 _18115_ (.A(_14323_),
    .B(_14236_),
    .Y(_14356_));
 sky130_fd_sc_hd__o21ai_1 _18116_ (.A1(_14354_),
    .A2(_14355_),
    .B1(_14356_),
    .Y(_03045_));
 sky130_fd_sc_hd__clkbuf_4 _18117_ (.A(\pcpi_mul.rs1[17] ),
    .X(_14357_));
 sky130_fd_sc_hd__clkinv_4 _18118_ (.A(_14357_),
    .Y(_14358_));
 sky130_fd_sc_hd__buf_4 _18119_ (.A(_14358_),
    .X(_14359_));
 sky130_fd_sc_hd__buf_6 _18120_ (.A(_14359_),
    .X(_14360_));
 sky130_fd_sc_hd__buf_6 _18121_ (.A(_14360_),
    .X(_14361_));
 sky130_fd_sc_hd__clkbuf_2 _18122_ (.A(_12795_),
    .X(_14362_));
 sky130_fd_sc_hd__nand2_1 _18123_ (.A(_14362_),
    .B(_14238_),
    .Y(_14363_));
 sky130_fd_sc_hd__o21ai_1 _18124_ (.A1(_14361_),
    .A2(_14355_),
    .B1(_14363_),
    .Y(_03044_));
 sky130_vsdinv _18125_ (.A(\pcpi_mul.rs1[16] ),
    .Y(_14364_));
 sky130_fd_sc_hd__buf_2 _18126_ (.A(_14364_),
    .X(_14365_));
 sky130_fd_sc_hd__buf_4 _18127_ (.A(_14365_),
    .X(_14366_));
 sky130_fd_sc_hd__buf_6 _18128_ (.A(_14366_),
    .X(_14367_));
 sky130_fd_sc_hd__buf_6 _18129_ (.A(_14367_),
    .X(_14368_));
 sky130_fd_sc_hd__nand2_1 _18130_ (.A(_14362_),
    .B(_14240_),
    .Y(_14369_));
 sky130_fd_sc_hd__o21ai_1 _18131_ (.A1(_14368_),
    .A2(_14355_),
    .B1(_14369_),
    .Y(_03043_));
 sky130_fd_sc_hd__clkbuf_2 _18132_ (.A(\pcpi_mul.rs1[15] ),
    .X(_14370_));
 sky130_vsdinv _18133_ (.A(_14370_),
    .Y(_14371_));
 sky130_fd_sc_hd__buf_4 _18134_ (.A(_14371_),
    .X(_14372_));
 sky130_fd_sc_hd__buf_4 _18135_ (.A(_14372_),
    .X(_14373_));
 sky130_fd_sc_hd__buf_6 _18136_ (.A(_14373_),
    .X(_14374_));
 sky130_fd_sc_hd__nand2_1 _18137_ (.A(_14362_),
    .B(_14241_),
    .Y(_14375_));
 sky130_fd_sc_hd__o21ai_1 _18138_ (.A1(_14374_),
    .A2(_14355_),
    .B1(_14375_),
    .Y(_03042_));
 sky130_fd_sc_hd__buf_2 _18139_ (.A(\pcpi_mul.rs1[14] ),
    .X(_14376_));
 sky130_vsdinv _18140_ (.A(_14376_),
    .Y(_14377_));
 sky130_fd_sc_hd__buf_4 _18141_ (.A(_14377_),
    .X(_14378_));
 sky130_fd_sc_hd__buf_6 _18142_ (.A(_14378_),
    .X(_14379_));
 sky130_fd_sc_hd__nand2_1 _18143_ (.A(_14362_),
    .B(_14242_),
    .Y(_14380_));
 sky130_fd_sc_hd__o21ai_1 _18144_ (.A1(_14379_),
    .A2(_14355_),
    .B1(_14380_),
    .Y(_03041_));
 sky130_fd_sc_hd__buf_2 _18145_ (.A(\pcpi_mul.rs1[13] ),
    .X(_14381_));
 sky130_vsdinv _18146_ (.A(_14381_),
    .Y(_14382_));
 sky130_fd_sc_hd__clkbuf_4 _18147_ (.A(_14382_),
    .X(_14383_));
 sky130_fd_sc_hd__buf_4 _18148_ (.A(_14383_),
    .X(_14384_));
 sky130_fd_sc_hd__clkbuf_8 _18149_ (.A(_14384_),
    .X(_14385_));
 sky130_fd_sc_hd__nand2_1 _18150_ (.A(_14362_),
    .B(_14243_),
    .Y(_14386_));
 sky130_fd_sc_hd__o21ai_1 _18151_ (.A1(_14385_),
    .A2(_14355_),
    .B1(_14386_),
    .Y(_03040_));
 sky130_fd_sc_hd__clkbuf_4 _18152_ (.A(\pcpi_mul.rs1[12] ),
    .X(_14387_));
 sky130_vsdinv _18153_ (.A(_14387_),
    .Y(_14388_));
 sky130_fd_sc_hd__buf_4 _18154_ (.A(_14388_),
    .X(_14389_));
 sky130_fd_sc_hd__buf_6 _18155_ (.A(_14389_),
    .X(_14390_));
 sky130_fd_sc_hd__clkbuf_2 _18156_ (.A(_14078_),
    .X(_14391_));
 sky130_fd_sc_hd__nand2_1 _18157_ (.A(_14362_),
    .B(_14245_),
    .Y(_14392_));
 sky130_fd_sc_hd__o21ai_1 _18158_ (.A1(_14390_),
    .A2(_14391_),
    .B1(_14392_),
    .Y(_03039_));
 sky130_vsdinv _18159_ (.A(\pcpi_mul.rs1[11] ),
    .Y(_14393_));
 sky130_fd_sc_hd__buf_4 _18160_ (.A(_14393_),
    .X(_14394_));
 sky130_fd_sc_hd__buf_4 _18161_ (.A(_14394_),
    .X(_14395_));
 sky130_fd_sc_hd__clkbuf_2 _18162_ (.A(_12795_),
    .X(_14396_));
 sky130_fd_sc_hd__nand2_1 _18163_ (.A(_14396_),
    .B(_14246_),
    .Y(_14397_));
 sky130_fd_sc_hd__o21ai_1 _18164_ (.A1(_14395_),
    .A2(_14391_),
    .B1(_14397_),
    .Y(_03038_));
 sky130_fd_sc_hd__clkbuf_2 _18165_ (.A(\pcpi_mul.rs1[10] ),
    .X(_14398_));
 sky130_fd_sc_hd__inv_2 _18166_ (.A(_14398_),
    .Y(_14399_));
 sky130_fd_sc_hd__clkbuf_4 _18167_ (.A(_14399_),
    .X(_14400_));
 sky130_fd_sc_hd__buf_4 _18168_ (.A(_14400_),
    .X(_14401_));
 sky130_fd_sc_hd__nand2_1 _18169_ (.A(_14396_),
    .B(_14247_),
    .Y(_14402_));
 sky130_fd_sc_hd__o21ai_1 _18170_ (.A1(_14401_),
    .A2(_14391_),
    .B1(_14402_),
    .Y(_03037_));
 sky130_vsdinv _18171_ (.A(\pcpi_mul.rs1[9] ),
    .Y(_14403_));
 sky130_fd_sc_hd__clkbuf_2 _18172_ (.A(_14403_),
    .X(_14404_));
 sky130_fd_sc_hd__buf_4 _18173_ (.A(_14404_),
    .X(_14405_));
 sky130_fd_sc_hd__buf_6 _18174_ (.A(_14405_),
    .X(_14406_));
 sky130_fd_sc_hd__nand2_1 _18175_ (.A(_14396_),
    .B(_14249_),
    .Y(_14407_));
 sky130_fd_sc_hd__o21ai_1 _18176_ (.A1(_14406_),
    .A2(_14391_),
    .B1(_14407_),
    .Y(_03036_));
 sky130_fd_sc_hd__clkbuf_2 _18177_ (.A(\pcpi_mul.rs1[8] ),
    .X(_14408_));
 sky130_vsdinv _18178_ (.A(_14408_),
    .Y(_14409_));
 sky130_fd_sc_hd__buf_2 _18179_ (.A(_14409_),
    .X(_14410_));
 sky130_fd_sc_hd__buf_4 _18180_ (.A(_14410_),
    .X(_14411_));
 sky130_fd_sc_hd__buf_6 _18181_ (.A(_14411_),
    .X(_14412_));
 sky130_fd_sc_hd__nand2_1 _18182_ (.A(_14396_),
    .B(_14251_),
    .Y(_14413_));
 sky130_fd_sc_hd__o21ai_1 _18183_ (.A1(_14412_),
    .A2(_14391_),
    .B1(_14413_),
    .Y(_03035_));
 sky130_fd_sc_hd__clkbuf_4 _18184_ (.A(\pcpi_mul.rs1[7] ),
    .X(_14414_));
 sky130_vsdinv _18185_ (.A(_14414_),
    .Y(_14415_));
 sky130_fd_sc_hd__buf_2 _18186_ (.A(_14415_),
    .X(_14416_));
 sky130_fd_sc_hd__clkbuf_4 _18187_ (.A(_14416_),
    .X(_14417_));
 sky130_fd_sc_hd__buf_6 _18188_ (.A(_14417_),
    .X(_14418_));
 sky130_fd_sc_hd__nand2_1 _18189_ (.A(_14396_),
    .B(_14253_),
    .Y(_14419_));
 sky130_fd_sc_hd__o21ai_1 _18190_ (.A1(_14418_),
    .A2(_14391_),
    .B1(_14419_),
    .Y(_03034_));
 sky130_fd_sc_hd__clkbuf_2 _18191_ (.A(\pcpi_mul.rs1[6] ),
    .X(_14420_));
 sky130_vsdinv _18192_ (.A(_14420_),
    .Y(_14421_));
 sky130_fd_sc_hd__clkbuf_4 _18193_ (.A(_14421_),
    .X(_14422_));
 sky130_fd_sc_hd__buf_6 _18194_ (.A(_14422_),
    .X(_14423_));
 sky130_fd_sc_hd__buf_2 _18195_ (.A(_14078_),
    .X(_14424_));
 sky130_fd_sc_hd__nand2_2 _18196_ (.A(_14396_),
    .B(_14256_),
    .Y(_14425_));
 sky130_fd_sc_hd__o21ai_1 _18197_ (.A1(_14423_),
    .A2(_14424_),
    .B1(_14425_),
    .Y(_03033_));
 sky130_fd_sc_hd__buf_2 _18198_ (.A(\pcpi_mul.rs1[5] ),
    .X(_14426_));
 sky130_vsdinv _18199_ (.A(_14426_),
    .Y(_14427_));
 sky130_fd_sc_hd__clkbuf_4 _18200_ (.A(_14427_),
    .X(_14428_));
 sky130_fd_sc_hd__buf_6 _18201_ (.A(_14428_),
    .X(_14429_));
 sky130_fd_sc_hd__clkbuf_4 _18202_ (.A(_12795_),
    .X(_14430_));
 sky130_fd_sc_hd__nand2_1 _18203_ (.A(_14430_),
    .B(_14257_),
    .Y(_14431_));
 sky130_fd_sc_hd__o21ai_1 _18204_ (.A1(_14429_),
    .A2(_14424_),
    .B1(_14431_),
    .Y(_03032_));
 sky130_fd_sc_hd__clkbuf_4 _18205_ (.A(\pcpi_mul.rs1[4] ),
    .X(_14432_));
 sky130_vsdinv _18206_ (.A(_14432_),
    .Y(_14433_));
 sky130_fd_sc_hd__clkbuf_4 _18207_ (.A(_14433_),
    .X(_14434_));
 sky130_fd_sc_hd__buf_6 _18208_ (.A(_14434_),
    .X(_14435_));
 sky130_fd_sc_hd__nand2_2 _18209_ (.A(_14430_),
    .B(_14259_),
    .Y(_14436_));
 sky130_fd_sc_hd__o21ai_1 _18210_ (.A1(_14435_),
    .A2(_14424_),
    .B1(_14436_),
    .Y(_03031_));
 sky130_vsdinv _18211_ (.A(\pcpi_mul.rs1[3] ),
    .Y(_14437_));
 sky130_fd_sc_hd__clkbuf_4 _18212_ (.A(_14437_),
    .X(_14438_));
 sky130_fd_sc_hd__buf_4 _18213_ (.A(_14438_),
    .X(_14439_));
 sky130_fd_sc_hd__nand2_2 _18214_ (.A(_14430_),
    .B(_14260_),
    .Y(_14440_));
 sky130_fd_sc_hd__o21ai_1 _18215_ (.A1(_14439_),
    .A2(_14424_),
    .B1(_14440_),
    .Y(_03030_));
 sky130_fd_sc_hd__buf_2 _18216_ (.A(\pcpi_mul.rs1[2] ),
    .X(_14441_));
 sky130_vsdinv _18217_ (.A(_14441_),
    .Y(_14442_));
 sky130_fd_sc_hd__buf_4 _18218_ (.A(_14442_),
    .X(_14443_));
 sky130_fd_sc_hd__buf_6 _18219_ (.A(_14443_),
    .X(_14444_));
 sky130_fd_sc_hd__buf_4 _18220_ (.A(_14444_),
    .X(_14445_));
 sky130_fd_sc_hd__nand2_2 _18221_ (.A(_14430_),
    .B(_14262_),
    .Y(_14446_));
 sky130_fd_sc_hd__o21ai_1 _18222_ (.A1(_14445_),
    .A2(_14424_),
    .B1(_14446_),
    .Y(_03029_));
 sky130_fd_sc_hd__buf_4 _18223_ (.A(\pcpi_mul.rs1[1] ),
    .X(_14447_));
 sky130_fd_sc_hd__buf_2 _18224_ (.A(_14447_),
    .X(_14448_));
 sky130_vsdinv _18225_ (.A(_14448_),
    .Y(_14449_));
 sky130_fd_sc_hd__nand2_1 _18226_ (.A(_14430_),
    .B(_14265_),
    .Y(_14450_));
 sky130_fd_sc_hd__o21ai_1 _18227_ (.A1(_14449_),
    .A2(_14424_),
    .B1(_14450_),
    .Y(_03028_));
 sky130_vsdinv _18228_ (.A(\pcpi_mul.rs1[0] ),
    .Y(_14451_));
 sky130_fd_sc_hd__buf_4 _18229_ (.A(_14451_),
    .X(_14452_));
 sky130_fd_sc_hd__buf_4 _18230_ (.A(_14452_),
    .X(_14453_));
 sky130_fd_sc_hd__buf_6 _18231_ (.A(_14453_),
    .X(_14454_));
 sky130_fd_sc_hd__nand2_1 _18232_ (.A(_14430_),
    .B(_14269_),
    .Y(_14455_));
 sky130_fd_sc_hd__o21ai_1 _18233_ (.A1(_14454_),
    .A2(_12794_),
    .B1(_14455_),
    .Y(_03027_));
 sky130_fd_sc_hd__clkbuf_2 _18234_ (.A(\cpuregs_wrdata[31] ),
    .X(_14456_));
 sky130_fd_sc_hd__nand2_1 _18235_ (.A(_13786_),
    .B(_13746_),
    .Y(_14457_));
 sky130_fd_sc_hd__buf_8 _18236_ (.A(_14457_),
    .X(_14458_));
 sky130_fd_sc_hd__buf_4 _18237_ (.A(_14458_),
    .X(_14459_));
 sky130_fd_sc_hd__mux2_1 _18238_ (.A0(_14456_),
    .A1(\cpuregs[5][31] ),
    .S(_14459_),
    .X(_03026_));
 sky130_fd_sc_hd__clkbuf_2 _18239_ (.A(\cpuregs_wrdata[30] ),
    .X(_14460_));
 sky130_fd_sc_hd__mux2_1 _18240_ (.A0(_14460_),
    .A1(\cpuregs[5][30] ),
    .S(_14459_),
    .X(_03025_));
 sky130_fd_sc_hd__clkbuf_2 _18241_ (.A(\cpuregs_wrdata[29] ),
    .X(_14461_));
 sky130_fd_sc_hd__mux2_1 _18242_ (.A0(_14461_),
    .A1(\cpuregs[5][29] ),
    .S(_14459_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_2 _18243_ (.A(\cpuregs_wrdata[28] ),
    .X(_14462_));
 sky130_fd_sc_hd__mux2_1 _18244_ (.A0(_14462_),
    .A1(\cpuregs[5][28] ),
    .S(_14459_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_2 _18245_ (.A(\cpuregs_wrdata[27] ),
    .X(_14463_));
 sky130_fd_sc_hd__mux2_1 _18246_ (.A0(_14463_),
    .A1(\cpuregs[5][27] ),
    .S(_14459_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_2 _18247_ (.A(\cpuregs_wrdata[26] ),
    .X(_14464_));
 sky130_fd_sc_hd__mux2_1 _18248_ (.A0(_14464_),
    .A1(\cpuregs[5][26] ),
    .S(_14459_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_2 _18249_ (.A(\cpuregs_wrdata[25] ),
    .X(_14465_));
 sky130_fd_sc_hd__buf_2 _18250_ (.A(_14458_),
    .X(_14466_));
 sky130_fd_sc_hd__mux2_1 _18251_ (.A0(_14465_),
    .A1(\cpuregs[5][25] ),
    .S(_14466_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_2 _18252_ (.A(\cpuregs_wrdata[24] ),
    .X(_14467_));
 sky130_fd_sc_hd__mux2_1 _18253_ (.A0(_14467_),
    .A1(\cpuregs[5][24] ),
    .S(_14466_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_2 _18254_ (.A(\cpuregs_wrdata[23] ),
    .X(_14468_));
 sky130_fd_sc_hd__mux2_1 _18255_ (.A0(_14468_),
    .A1(\cpuregs[5][23] ),
    .S(_14466_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_2 _18256_ (.A(\cpuregs_wrdata[22] ),
    .X(_14469_));
 sky130_fd_sc_hd__mux2_1 _18257_ (.A0(_14469_),
    .A1(\cpuregs[5][22] ),
    .S(_14466_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_2 _18258_ (.A(\cpuregs_wrdata[21] ),
    .X(_14470_));
 sky130_fd_sc_hd__mux2_1 _18259_ (.A0(_14470_),
    .A1(\cpuregs[5][21] ),
    .S(_14466_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_2 _18260_ (.A(\cpuregs_wrdata[20] ),
    .X(_14471_));
 sky130_fd_sc_hd__mux2_1 _18261_ (.A0(_14471_),
    .A1(\cpuregs[5][20] ),
    .S(_14466_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_2 _18262_ (.A(\cpuregs_wrdata[19] ),
    .X(_14472_));
 sky130_fd_sc_hd__buf_2 _18263_ (.A(_14458_),
    .X(_14473_));
 sky130_fd_sc_hd__mux2_1 _18264_ (.A0(_14472_),
    .A1(\cpuregs[5][19] ),
    .S(_14473_),
    .X(_03014_));
 sky130_fd_sc_hd__buf_2 _18265_ (.A(\cpuregs_wrdata[18] ),
    .X(_14474_));
 sky130_fd_sc_hd__mux2_1 _18266_ (.A0(_14474_),
    .A1(\cpuregs[5][18] ),
    .S(_14473_),
    .X(_03013_));
 sky130_fd_sc_hd__buf_2 _18267_ (.A(\cpuregs_wrdata[17] ),
    .X(_14475_));
 sky130_fd_sc_hd__mux2_1 _18268_ (.A0(_14475_),
    .A1(\cpuregs[5][17] ),
    .S(_14473_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_2 _18269_ (.A(\cpuregs_wrdata[16] ),
    .X(_14476_));
 sky130_fd_sc_hd__mux2_1 _18270_ (.A0(_14476_),
    .A1(\cpuregs[5][16] ),
    .S(_14473_),
    .X(_03011_));
 sky130_fd_sc_hd__clkbuf_2 _18271_ (.A(\cpuregs_wrdata[15] ),
    .X(_14477_));
 sky130_fd_sc_hd__mux2_1 _18272_ (.A0(_14477_),
    .A1(\cpuregs[5][15] ),
    .S(_14473_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_2 _18273_ (.A(\cpuregs_wrdata[14] ),
    .X(_14478_));
 sky130_fd_sc_hd__mux2_1 _18274_ (.A0(_14478_),
    .A1(\cpuregs[5][14] ),
    .S(_14473_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_2 _18275_ (.A(\cpuregs_wrdata[13] ),
    .X(_14479_));
 sky130_fd_sc_hd__buf_4 _18276_ (.A(_14458_),
    .X(_14480_));
 sky130_fd_sc_hd__mux2_1 _18277_ (.A0(_14479_),
    .A1(\cpuregs[5][13] ),
    .S(_14480_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_2 _18278_ (.A(\cpuregs_wrdata[12] ),
    .X(_14481_));
 sky130_fd_sc_hd__mux2_1 _18279_ (.A0(_14481_),
    .A1(\cpuregs[5][12] ),
    .S(_14480_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_2 _18280_ (.A(\cpuregs_wrdata[11] ),
    .X(_14482_));
 sky130_fd_sc_hd__mux2_1 _18281_ (.A0(_14482_),
    .A1(\cpuregs[5][11] ),
    .S(_14480_),
    .X(_03006_));
 sky130_fd_sc_hd__clkbuf_2 _18282_ (.A(\cpuregs_wrdata[10] ),
    .X(_14483_));
 sky130_fd_sc_hd__mux2_1 _18283_ (.A0(_14483_),
    .A1(\cpuregs[5][10] ),
    .S(_14480_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_2 _18284_ (.A(\cpuregs_wrdata[9] ),
    .X(_14484_));
 sky130_fd_sc_hd__mux2_1 _18285_ (.A0(_14484_),
    .A1(\cpuregs[5][9] ),
    .S(_14480_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_2 _18286_ (.A(\cpuregs_wrdata[8] ),
    .X(_14485_));
 sky130_fd_sc_hd__mux2_1 _18287_ (.A0(_14485_),
    .A1(\cpuregs[5][8] ),
    .S(_14480_),
    .X(_03003_));
 sky130_fd_sc_hd__clkbuf_2 _18288_ (.A(\cpuregs_wrdata[7] ),
    .X(_14486_));
 sky130_fd_sc_hd__clkbuf_4 _18289_ (.A(_14457_),
    .X(_14487_));
 sky130_fd_sc_hd__mux2_1 _18290_ (.A0(_14486_),
    .A1(\cpuregs[5][7] ),
    .S(_14487_),
    .X(_03002_));
 sky130_fd_sc_hd__clkbuf_2 _18291_ (.A(\cpuregs_wrdata[6] ),
    .X(_14488_));
 sky130_fd_sc_hd__mux2_1 _18292_ (.A0(_14488_),
    .A1(\cpuregs[5][6] ),
    .S(_14487_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_2 _18293_ (.A(\cpuregs_wrdata[5] ),
    .X(_14489_));
 sky130_fd_sc_hd__mux2_1 _18294_ (.A0(_14489_),
    .A1(\cpuregs[5][5] ),
    .S(_14487_),
    .X(_03000_));
 sky130_fd_sc_hd__clkbuf_2 _18295_ (.A(\cpuregs_wrdata[4] ),
    .X(_14490_));
 sky130_fd_sc_hd__mux2_1 _18296_ (.A0(_14490_),
    .A1(\cpuregs[5][4] ),
    .S(_14487_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_2 _18297_ (.A(\cpuregs_wrdata[3] ),
    .X(_14491_));
 sky130_fd_sc_hd__mux2_1 _18298_ (.A0(_14491_),
    .A1(\cpuregs[5][3] ),
    .S(_14487_),
    .X(_02998_));
 sky130_fd_sc_hd__clkbuf_2 _18299_ (.A(\cpuregs_wrdata[2] ),
    .X(_14492_));
 sky130_fd_sc_hd__mux2_1 _18300_ (.A0(_14492_),
    .A1(\cpuregs[5][2] ),
    .S(_14487_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_2 _18301_ (.A(\cpuregs_wrdata[1] ),
    .X(_14493_));
 sky130_fd_sc_hd__mux2_1 _18302_ (.A0(_14493_),
    .A1(\cpuregs[5][1] ),
    .S(_14458_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_2 _18303_ (.A(\cpuregs_wrdata[0] ),
    .X(_14494_));
 sky130_fd_sc_hd__mux2_1 _18304_ (.A0(_14494_),
    .A1(\cpuregs[5][0] ),
    .S(_14458_),
    .X(_02995_));
 sky130_fd_sc_hd__nand2_1 _18305_ (.A(_13743_),
    .B(_13738_),
    .Y(_14495_));
 sky130_fd_sc_hd__buf_6 _18306_ (.A(_14495_),
    .X(_14496_));
 sky130_fd_sc_hd__buf_4 _18307_ (.A(_14496_),
    .X(_14497_));
 sky130_fd_sc_hd__mux2_1 _18308_ (.A0(_14456_),
    .A1(\cpuregs[2][31] ),
    .S(_14497_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _18309_ (.A0(_14460_),
    .A1(\cpuregs[2][30] ),
    .S(_14497_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_1 _18310_ (.A0(_14461_),
    .A1(\cpuregs[2][29] ),
    .S(_14497_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_1 _18311_ (.A0(_14462_),
    .A1(\cpuregs[2][28] ),
    .S(_14497_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _18312_ (.A0(_14463_),
    .A1(\cpuregs[2][27] ),
    .S(_14497_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _18313_ (.A0(_14464_),
    .A1(\cpuregs[2][26] ),
    .S(_14497_),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_4 _18314_ (.A(_14496_),
    .X(_14498_));
 sky130_fd_sc_hd__mux2_1 _18315_ (.A0(_14465_),
    .A1(\cpuregs[2][25] ),
    .S(_14498_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _18316_ (.A0(_14467_),
    .A1(\cpuregs[2][24] ),
    .S(_14498_),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_1 _18317_ (.A0(_14468_),
    .A1(\cpuregs[2][23] ),
    .S(_14498_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _18318_ (.A0(_14469_),
    .A1(\cpuregs[2][22] ),
    .S(_14498_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_1 _18319_ (.A0(_14470_),
    .A1(\cpuregs[2][21] ),
    .S(_14498_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _18320_ (.A0(_14471_),
    .A1(\cpuregs[2][20] ),
    .S(_14498_),
    .X(_02983_));
 sky130_fd_sc_hd__clkbuf_4 _18321_ (.A(_14496_),
    .X(_14499_));
 sky130_fd_sc_hd__mux2_1 _18322_ (.A0(_14472_),
    .A1(\cpuregs[2][19] ),
    .S(_14499_),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_1 _18323_ (.A0(_14474_),
    .A1(\cpuregs[2][18] ),
    .S(_14499_),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_1 _18324_ (.A0(_14475_),
    .A1(\cpuregs[2][17] ),
    .S(_14499_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _18325_ (.A0(_14476_),
    .A1(\cpuregs[2][16] ),
    .S(_14499_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _18326_ (.A0(_14477_),
    .A1(\cpuregs[2][15] ),
    .S(_14499_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_1 _18327_ (.A0(_14478_),
    .A1(\cpuregs[2][14] ),
    .S(_14499_),
    .X(_02977_));
 sky130_fd_sc_hd__clkbuf_4 _18328_ (.A(_14496_),
    .X(_14500_));
 sky130_fd_sc_hd__mux2_1 _18329_ (.A0(_14479_),
    .A1(\cpuregs[2][13] ),
    .S(_14500_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _18330_ (.A0(_14481_),
    .A1(\cpuregs[2][12] ),
    .S(_14500_),
    .X(_02975_));
 sky130_fd_sc_hd__mux2_1 _18331_ (.A0(_14482_),
    .A1(\cpuregs[2][11] ),
    .S(_14500_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_1 _18332_ (.A0(_14483_),
    .A1(\cpuregs[2][10] ),
    .S(_14500_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _18333_ (.A0(_14484_),
    .A1(\cpuregs[2][9] ),
    .S(_14500_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _18334_ (.A0(_14485_),
    .A1(\cpuregs[2][8] ),
    .S(_14500_),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_4 _18335_ (.A(_14495_),
    .X(_14501_));
 sky130_fd_sc_hd__mux2_1 _18336_ (.A0(_14486_),
    .A1(\cpuregs[2][7] ),
    .S(_14501_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _18337_ (.A0(_14488_),
    .A1(\cpuregs[2][6] ),
    .S(_14501_),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _18338_ (.A0(_14489_),
    .A1(\cpuregs[2][5] ),
    .S(_14501_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _18339_ (.A0(_14490_),
    .A1(\cpuregs[2][4] ),
    .S(_14501_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _18340_ (.A0(_14491_),
    .A1(\cpuregs[2][3] ),
    .S(_14501_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_1 _18341_ (.A0(_14492_),
    .A1(\cpuregs[2][2] ),
    .S(_14501_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _18342_ (.A0(_14493_),
    .A1(\cpuregs[2][1] ),
    .S(_14496_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _18343_ (.A0(_14494_),
    .A1(\cpuregs[2][0] ),
    .S(_14496_),
    .X(_02963_));
 sky130_fd_sc_hd__clkbuf_2 _18344_ (.A(_12629_),
    .X(_14502_));
 sky130_fd_sc_hd__clkbuf_2 _18345_ (.A(_14502_),
    .X(mem_xfer));
 sky130_fd_sc_hd__mux2_1 _18346_ (.A0(_14207_),
    .A1(net57),
    .S(net444),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _18347_ (.A0(\mem_rdata_q[30] ),
    .A1(net497),
    .S(net445),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _18348_ (.A0(_13014_),
    .A1(net54),
    .S(net445),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _18349_ (.A0(\mem_rdata_q[28] ),
    .A1(net53),
    .S(net444),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_1 _18350_ (.A0(_14141_),
    .A1(net52),
    .S(net444),
    .X(_02958_));
 sky130_fd_sc_hd__buf_2 _18351_ (.A(_14502_),
    .X(_14503_));
 sky130_fd_sc_hd__mux2_1 _18352_ (.A0(\mem_rdata_q[26] ),
    .A1(net51),
    .S(_14503_),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_1 _18353_ (.A0(_14154_),
    .A1(net50),
    .S(_14503_),
    .X(_02956_));
 sky130_fd_sc_hd__mux2_1 _18354_ (.A0(\mem_rdata_q[24] ),
    .A1(net49),
    .S(_14503_),
    .X(_02955_));
 sky130_fd_sc_hd__mux2_1 _18355_ (.A0(\mem_rdata_q[23] ),
    .A1(net48),
    .S(_14503_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _18356_ (.A0(\mem_rdata_q[22] ),
    .A1(net47),
    .S(_14503_),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_1 _18357_ (.A0(\mem_rdata_q[21] ),
    .A1(net46),
    .S(_14503_),
    .X(_02952_));
 sky130_fd_sc_hd__buf_2 _18358_ (.A(_14502_),
    .X(_14504_));
 sky130_fd_sc_hd__mux2_1 _18359_ (.A0(\mem_rdata_q[20] ),
    .A1(net45),
    .S(_14504_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _18360_ (.A0(\mem_rdata_q[19] ),
    .A1(net498),
    .S(_14504_),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_1 _18361_ (.A0(\mem_rdata_q[18] ),
    .A1(net42),
    .S(_14504_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _18362_ (.A0(\mem_rdata_q[17] ),
    .A1(net499),
    .S(_14504_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _18363_ (.A0(\mem_rdata_q[16] ),
    .A1(net40),
    .S(_14504_),
    .X(_02947_));
 sky130_fd_sc_hd__mux2_1 _18364_ (.A0(\mem_rdata_q[15] ),
    .A1(net500),
    .S(_14504_),
    .X(_02946_));
 sky130_fd_sc_hd__buf_2 _18365_ (.A(_12629_),
    .X(_14505_));
 sky130_fd_sc_hd__mux2_1 _18366_ (.A0(_12990_),
    .A1(net38),
    .S(_14505_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_1 _18367_ (.A0(_12992_),
    .A1(net37),
    .S(_14505_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _18368_ (.A0(_12994_),
    .A1(net36),
    .S(_14505_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _18369_ (.A0(\mem_rdata_q[11] ),
    .A1(net35),
    .S(_14505_),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_1 _18370_ (.A0(\mem_rdata_q[10] ),
    .A1(net34),
    .S(_14505_),
    .X(_02941_));
 sky130_fd_sc_hd__mux2_1 _18371_ (.A0(\mem_rdata_q[9] ),
    .A1(net64),
    .S(_14505_),
    .X(_02940_));
 sky130_fd_sc_hd__buf_2 _18372_ (.A(_12629_),
    .X(_14506_));
 sky130_fd_sc_hd__mux2_1 _18373_ (.A0(\mem_rdata_q[8] ),
    .A1(net63),
    .S(_14506_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _18374_ (.A0(\mem_rdata_q[7] ),
    .A1(net62),
    .S(_14506_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _18375_ (.A0(\mem_rdata_q[6] ),
    .A1(net61),
    .S(_14506_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _18376_ (.A0(\mem_rdata_q[5] ),
    .A1(net60),
    .S(_14506_),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_1 _18377_ (.A0(\mem_rdata_q[4] ),
    .A1(net59),
    .S(_14506_),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_1 _18378_ (.A0(\mem_rdata_q[3] ),
    .A1(net58),
    .S(_14506_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_1 _18379_ (.A0(\mem_rdata_q[2] ),
    .A1(net55),
    .S(_14502_),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_1 _18380_ (.A0(\mem_rdata_q[1] ),
    .A1(net44),
    .S(_14502_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _18381_ (.A0(\mem_rdata_q[0] ),
    .A1(net33),
    .S(_14502_),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_1 _18382_ (.A(_13743_),
    .B(_13849_),
    .Y(_14507_));
 sky130_fd_sc_hd__buf_6 _18383_ (.A(_14507_),
    .X(_14508_));
 sky130_fd_sc_hd__clkbuf_4 _18384_ (.A(_14508_),
    .X(_14509_));
 sky130_fd_sc_hd__mux2_1 _18385_ (.A0(_14456_),
    .A1(\cpuregs[18][31] ),
    .S(_14509_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _18386_ (.A0(_14460_),
    .A1(\cpuregs[18][30] ),
    .S(_14509_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_1 _18387_ (.A0(_14461_),
    .A1(\cpuregs[18][29] ),
    .S(_14509_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_1 _18388_ (.A0(_14462_),
    .A1(\cpuregs[18][28] ),
    .S(_14509_),
    .X(_02927_));
 sky130_fd_sc_hd__mux2_1 _18389_ (.A0(_14463_),
    .A1(\cpuregs[18][27] ),
    .S(_14509_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _18390_ (.A0(_14464_),
    .A1(\cpuregs[18][26] ),
    .S(_14509_),
    .X(_02925_));
 sky130_fd_sc_hd__clkbuf_4 _18391_ (.A(_14508_),
    .X(_14510_));
 sky130_fd_sc_hd__mux2_1 _18392_ (.A0(_14465_),
    .A1(\cpuregs[18][25] ),
    .S(_14510_),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_1 _18393_ (.A0(_14467_),
    .A1(\cpuregs[18][24] ),
    .S(_14510_),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _18394_ (.A0(_14468_),
    .A1(\cpuregs[18][23] ),
    .S(_14510_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _18395_ (.A0(_14469_),
    .A1(\cpuregs[18][22] ),
    .S(_14510_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _18396_ (.A0(_14470_),
    .A1(\cpuregs[18][21] ),
    .S(_14510_),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_1 _18397_ (.A0(_14471_),
    .A1(\cpuregs[18][20] ),
    .S(_14510_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_4 _18398_ (.A(_14508_),
    .X(_14511_));
 sky130_fd_sc_hd__mux2_1 _18399_ (.A0(_14472_),
    .A1(\cpuregs[18][19] ),
    .S(_14511_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _18400_ (.A0(_14474_),
    .A1(\cpuregs[18][18] ),
    .S(_14511_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _18401_ (.A0(_14475_),
    .A1(\cpuregs[18][17] ),
    .S(_14511_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _18402_ (.A0(_14476_),
    .A1(\cpuregs[18][16] ),
    .S(_14511_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _18403_ (.A0(_14477_),
    .A1(\cpuregs[18][15] ),
    .S(_14511_),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _18404_ (.A0(_14478_),
    .A1(\cpuregs[18][14] ),
    .S(_14511_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_4 _18405_ (.A(_14508_),
    .X(_14512_));
 sky130_fd_sc_hd__mux2_1 _18406_ (.A0(_14479_),
    .A1(\cpuregs[18][13] ),
    .S(_14512_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _18407_ (.A0(_14481_),
    .A1(\cpuregs[18][12] ),
    .S(_14512_),
    .X(_02911_));
 sky130_fd_sc_hd__mux2_1 _18408_ (.A0(_14482_),
    .A1(\cpuregs[18][11] ),
    .S(_14512_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _18409_ (.A0(_14483_),
    .A1(\cpuregs[18][10] ),
    .S(_14512_),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_1 _18410_ (.A0(_14484_),
    .A1(\cpuregs[18][9] ),
    .S(_14512_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _18411_ (.A0(_14485_),
    .A1(\cpuregs[18][8] ),
    .S(_14512_),
    .X(_02907_));
 sky130_fd_sc_hd__clkbuf_4 _18412_ (.A(_14507_),
    .X(_14513_));
 sky130_fd_sc_hd__mux2_1 _18413_ (.A0(_14486_),
    .A1(\cpuregs[18][7] ),
    .S(_14513_),
    .X(_02906_));
 sky130_fd_sc_hd__mux2_1 _18414_ (.A0(_14488_),
    .A1(\cpuregs[18][6] ),
    .S(_14513_),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_1 _18415_ (.A0(_14489_),
    .A1(\cpuregs[18][5] ),
    .S(_14513_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _18416_ (.A0(_14490_),
    .A1(\cpuregs[18][4] ),
    .S(_14513_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _18417_ (.A0(_14491_),
    .A1(\cpuregs[18][3] ),
    .S(_14513_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_1 _18418_ (.A0(_14492_),
    .A1(\cpuregs[18][2] ),
    .S(_14513_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _18419_ (.A0(_14493_),
    .A1(\cpuregs[18][1] ),
    .S(_14508_),
    .X(_02900_));
 sky130_fd_sc_hd__mux2_1 _18420_ (.A0(_14494_),
    .A1(\cpuregs[18][0] ),
    .S(_14508_),
    .X(_02899_));
 sky130_fd_sc_hd__nand2_1 _18421_ (.A(_13743_),
    .B(_13787_),
    .Y(_14514_));
 sky130_fd_sc_hd__buf_6 _18422_ (.A(_14514_),
    .X(_14515_));
 sky130_fd_sc_hd__clkbuf_4 _18423_ (.A(_14515_),
    .X(_14516_));
 sky130_fd_sc_hd__mux2_1 _18424_ (.A0(_14456_),
    .A1(\cpuregs[10][31] ),
    .S(_14516_),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_1 _18425_ (.A0(_14460_),
    .A1(\cpuregs[10][30] ),
    .S(_14516_),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_1 _18426_ (.A0(_14461_),
    .A1(\cpuregs[10][29] ),
    .S(_14516_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _18427_ (.A0(_14462_),
    .A1(\cpuregs[10][28] ),
    .S(_14516_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _18428_ (.A0(_14463_),
    .A1(\cpuregs[10][27] ),
    .S(_14516_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _18429_ (.A0(_14464_),
    .A1(\cpuregs[10][26] ),
    .S(_14516_),
    .X(_02893_));
 sky130_fd_sc_hd__clkbuf_4 _18430_ (.A(_14515_),
    .X(_14517_));
 sky130_fd_sc_hd__mux2_1 _18431_ (.A0(_14465_),
    .A1(\cpuregs[10][25] ),
    .S(_14517_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _18432_ (.A0(_14467_),
    .A1(\cpuregs[10][24] ),
    .S(_14517_),
    .X(_02891_));
 sky130_fd_sc_hd__mux2_1 _18433_ (.A0(_14468_),
    .A1(\cpuregs[10][23] ),
    .S(_14517_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_1 _18434_ (.A0(_14469_),
    .A1(\cpuregs[10][22] ),
    .S(_14517_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_1 _18435_ (.A0(_14470_),
    .A1(\cpuregs[10][21] ),
    .S(_14517_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _18436_ (.A0(_14471_),
    .A1(\cpuregs[10][20] ),
    .S(_14517_),
    .X(_02887_));
 sky130_fd_sc_hd__clkbuf_4 _18437_ (.A(_14515_),
    .X(_14518_));
 sky130_fd_sc_hd__mux2_1 _18438_ (.A0(_14472_),
    .A1(\cpuregs[10][19] ),
    .S(_14518_),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_1 _18439_ (.A0(_14474_),
    .A1(\cpuregs[10][18] ),
    .S(_14518_),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_1 _18440_ (.A0(_14475_),
    .A1(\cpuregs[10][17] ),
    .S(_14518_),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_1 _18441_ (.A0(_14476_),
    .A1(\cpuregs[10][16] ),
    .S(_14518_),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _18442_ (.A0(_14477_),
    .A1(\cpuregs[10][15] ),
    .S(_14518_),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _18443_ (.A0(_14478_),
    .A1(\cpuregs[10][14] ),
    .S(_14518_),
    .X(_02881_));
 sky130_fd_sc_hd__clkbuf_4 _18444_ (.A(_14515_),
    .X(_14519_));
 sky130_fd_sc_hd__mux2_1 _18445_ (.A0(_14479_),
    .A1(\cpuregs[10][13] ),
    .S(_14519_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _18446_ (.A0(_14481_),
    .A1(\cpuregs[10][12] ),
    .S(_14519_),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _18447_ (.A0(_14482_),
    .A1(\cpuregs[10][11] ),
    .S(_14519_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _18448_ (.A0(_14483_),
    .A1(\cpuregs[10][10] ),
    .S(_14519_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _18449_ (.A0(_14484_),
    .A1(\cpuregs[10][9] ),
    .S(_14519_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _18450_ (.A0(_14485_),
    .A1(\cpuregs[10][8] ),
    .S(_14519_),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_4 _18451_ (.A(_14514_),
    .X(_14520_));
 sky130_fd_sc_hd__mux2_1 _18452_ (.A0(_14486_),
    .A1(\cpuregs[10][7] ),
    .S(_14520_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _18453_ (.A0(_14488_),
    .A1(\cpuregs[10][6] ),
    .S(_14520_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _18454_ (.A0(_14489_),
    .A1(\cpuregs[10][5] ),
    .S(_14520_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _18455_ (.A0(_14490_),
    .A1(\cpuregs[10][4] ),
    .S(_14520_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _18456_ (.A0(_14491_),
    .A1(\cpuregs[10][3] ),
    .S(_14520_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _18457_ (.A0(_14492_),
    .A1(\cpuregs[10][2] ),
    .S(_14520_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_1 _18458_ (.A0(_14493_),
    .A1(\cpuregs[10][1] ),
    .S(_14515_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _18459_ (.A0(_14494_),
    .A1(\cpuregs[10][0] ),
    .S(_14515_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_1 _18460_ (.A(\cpuregs[0][31] ),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_1 _18461_ (.A(\cpuregs[0][30] ),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _18462_ (.A(\cpuregs[0][29] ),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _18463_ (.A(\cpuregs[0][28] ),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _18464_ (.A(\cpuregs[0][27] ),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_1 _18465_ (.A(\cpuregs[0][26] ),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_1 _18466_ (.A(\cpuregs[0][25] ),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _18467_ (.A(\cpuregs[0][24] ),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _18468_ (.A(\cpuregs[0][23] ),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_1 _18469_ (.A(\cpuregs[0][22] ),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _18470_ (.A(\cpuregs[0][21] ),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_1 _18471_ (.A(\cpuregs[0][20] ),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _18472_ (.A(\cpuregs[0][19] ),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _18473_ (.A(\cpuregs[0][18] ),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _18474_ (.A(\cpuregs[0][17] ),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _18475_ (.A(\cpuregs[0][16] ),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _18476_ (.A(\cpuregs[0][15] ),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _18477_ (.A(\cpuregs[0][14] ),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _18478_ (.A(\cpuregs[0][13] ),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _18479_ (.A(\cpuregs[0][12] ),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _18480_ (.A(\cpuregs[0][11] ),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_1 _18481_ (.A(\cpuregs[0][10] ),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _18482_ (.A(\cpuregs[0][9] ),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _18483_ (.A(\cpuregs[0][8] ),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _18484_ (.A(\cpuregs[0][7] ),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _18485_ (.A(\cpuregs[0][6] ),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _18486_ (.A(\cpuregs[0][5] ),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _18487_ (.A(\cpuregs[0][4] ),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _18488_ (.A(\cpuregs[0][3] ),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _18489_ (.A(\cpuregs[0][2] ),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _18490_ (.A(\cpuregs[0][1] ),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _18491_ (.A(\cpuregs[0][0] ),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_1 _18492_ (.A(_13743_),
    .B(_13878_),
    .Y(_14521_));
 sky130_fd_sc_hd__buf_6 _18493_ (.A(_14521_),
    .X(_14522_));
 sky130_fd_sc_hd__clkbuf_4 _18494_ (.A(_14522_),
    .X(_14523_));
 sky130_fd_sc_hd__mux2_1 _18495_ (.A0(_14456_),
    .A1(\cpuregs[14][31] ),
    .S(_14523_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _18496_ (.A0(_14460_),
    .A1(\cpuregs[14][30] ),
    .S(_14523_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _18497_ (.A0(_14461_),
    .A1(\cpuregs[14][29] ),
    .S(_14523_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _18498_ (.A0(_14462_),
    .A1(\cpuregs[14][28] ),
    .S(_14523_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _18499_ (.A0(_14463_),
    .A1(\cpuregs[14][27] ),
    .S(_14523_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _18500_ (.A0(_14464_),
    .A1(\cpuregs[14][26] ),
    .S(_14523_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_4 _18501_ (.A(_14522_),
    .X(_14524_));
 sky130_fd_sc_hd__mux2_1 _18502_ (.A0(_14465_),
    .A1(\cpuregs[14][25] ),
    .S(_14524_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _18503_ (.A0(_14467_),
    .A1(\cpuregs[14][24] ),
    .S(_14524_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _18504_ (.A0(_14468_),
    .A1(\cpuregs[14][23] ),
    .S(_14524_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _18505_ (.A0(_14469_),
    .A1(\cpuregs[14][22] ),
    .S(_14524_),
    .X(_02825_));
 sky130_fd_sc_hd__mux2_1 _18506_ (.A0(_14470_),
    .A1(\cpuregs[14][21] ),
    .S(_14524_),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_1 _18507_ (.A0(_14471_),
    .A1(\cpuregs[14][20] ),
    .S(_14524_),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_4 _18508_ (.A(_14522_),
    .X(_14525_));
 sky130_fd_sc_hd__mux2_1 _18509_ (.A0(_14472_),
    .A1(\cpuregs[14][19] ),
    .S(_14525_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _18510_ (.A0(_14474_),
    .A1(\cpuregs[14][18] ),
    .S(_14525_),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_1 _18511_ (.A0(_14475_),
    .A1(\cpuregs[14][17] ),
    .S(_14525_),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_1 _18512_ (.A0(_14476_),
    .A1(\cpuregs[14][16] ),
    .S(_14525_),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _18513_ (.A0(_14477_),
    .A1(\cpuregs[14][15] ),
    .S(_14525_),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _18514_ (.A0(_14478_),
    .A1(\cpuregs[14][14] ),
    .S(_14525_),
    .X(_02817_));
 sky130_fd_sc_hd__buf_4 _18515_ (.A(_14522_),
    .X(_14526_));
 sky130_fd_sc_hd__mux2_1 _18516_ (.A0(_14479_),
    .A1(\cpuregs[14][13] ),
    .S(_14526_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _18517_ (.A0(_14481_),
    .A1(\cpuregs[14][12] ),
    .S(_14526_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _18518_ (.A0(_14482_),
    .A1(\cpuregs[14][11] ),
    .S(_14526_),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _18519_ (.A0(_14483_),
    .A1(\cpuregs[14][10] ),
    .S(_14526_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _18520_ (.A0(_14484_),
    .A1(\cpuregs[14][9] ),
    .S(_14526_),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _18521_ (.A0(_14485_),
    .A1(\cpuregs[14][8] ),
    .S(_14526_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_4 _18522_ (.A(_14521_),
    .X(_14527_));
 sky130_fd_sc_hd__mux2_1 _18523_ (.A0(_14486_),
    .A1(\cpuregs[14][7] ),
    .S(_14527_),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _18524_ (.A0(_14488_),
    .A1(\cpuregs[14][6] ),
    .S(_14527_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _18525_ (.A0(_14489_),
    .A1(\cpuregs[14][5] ),
    .S(_14527_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _18526_ (.A0(_14490_),
    .A1(\cpuregs[14][4] ),
    .S(_14527_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _18527_ (.A0(_14491_),
    .A1(\cpuregs[14][3] ),
    .S(_14527_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _18528_ (.A0(_14492_),
    .A1(\cpuregs[14][2] ),
    .S(_14527_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _18529_ (.A0(_14493_),
    .A1(\cpuregs[14][1] ),
    .S(_14522_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _18530_ (.A0(_14494_),
    .A1(\cpuregs[14][0] ),
    .S(_14522_),
    .X(_02803_));
 sky130_fd_sc_hd__nand3b_2 _18531_ (.A_N(_13742_),
    .B(_13739_),
    .C(_13787_),
    .Y(_14528_));
 sky130_fd_sc_hd__clkbuf_8 _18532_ (.A(_14528_),
    .X(_14529_));
 sky130_fd_sc_hd__clkbuf_4 _18533_ (.A(_14529_),
    .X(_14530_));
 sky130_fd_sc_hd__mux2_1 _18534_ (.A0(_14456_),
    .A1(\cpuregs[8][31] ),
    .S(_14530_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _18535_ (.A0(_14460_),
    .A1(\cpuregs[8][30] ),
    .S(_14530_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _18536_ (.A0(_14461_),
    .A1(\cpuregs[8][29] ),
    .S(_14530_),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_1 _18537_ (.A0(_14462_),
    .A1(\cpuregs[8][28] ),
    .S(_14530_),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _18538_ (.A0(_14463_),
    .A1(\cpuregs[8][27] ),
    .S(_14530_),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_1 _18539_ (.A0(_14464_),
    .A1(\cpuregs[8][26] ),
    .S(_14530_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_4 _18540_ (.A(_14529_),
    .X(_14531_));
 sky130_fd_sc_hd__mux2_1 _18541_ (.A0(_14465_),
    .A1(\cpuregs[8][25] ),
    .S(_14531_),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_1 _18542_ (.A0(_14467_),
    .A1(\cpuregs[8][24] ),
    .S(_14531_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _18543_ (.A0(_14468_),
    .A1(\cpuregs[8][23] ),
    .S(_14531_),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_1 _18544_ (.A0(_14469_),
    .A1(\cpuregs[8][22] ),
    .S(_14531_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_1 _18545_ (.A0(_14470_),
    .A1(\cpuregs[8][21] ),
    .S(_14531_),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_1 _18546_ (.A0(_14471_),
    .A1(\cpuregs[8][20] ),
    .S(_14531_),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_4 _18547_ (.A(_14529_),
    .X(_14532_));
 sky130_fd_sc_hd__mux2_1 _18548_ (.A0(_14472_),
    .A1(\cpuregs[8][19] ),
    .S(_14532_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _18549_ (.A0(_14474_),
    .A1(\cpuregs[8][18] ),
    .S(_14532_),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_1 _18550_ (.A0(_14475_),
    .A1(\cpuregs[8][17] ),
    .S(_14532_),
    .X(_02788_));
 sky130_fd_sc_hd__mux2_1 _18551_ (.A0(_14476_),
    .A1(\cpuregs[8][16] ),
    .S(_14532_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _18552_ (.A0(_14477_),
    .A1(\cpuregs[8][15] ),
    .S(_14532_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _18553_ (.A0(_14478_),
    .A1(\cpuregs[8][14] ),
    .S(_14532_),
    .X(_02785_));
 sky130_fd_sc_hd__clkbuf_4 _18554_ (.A(_14529_),
    .X(_14533_));
 sky130_fd_sc_hd__mux2_1 _18555_ (.A0(_14479_),
    .A1(\cpuregs[8][13] ),
    .S(_14533_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _18556_ (.A0(_14481_),
    .A1(\cpuregs[8][12] ),
    .S(_14533_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _18557_ (.A0(_14482_),
    .A1(\cpuregs[8][11] ),
    .S(_14533_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _18558_ (.A0(_14483_),
    .A1(\cpuregs[8][10] ),
    .S(_14533_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _18559_ (.A0(_14484_),
    .A1(\cpuregs[8][9] ),
    .S(_14533_),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_1 _18560_ (.A0(_14485_),
    .A1(\cpuregs[8][8] ),
    .S(_14533_),
    .X(_02779_));
 sky130_fd_sc_hd__clkbuf_4 _18561_ (.A(_14528_),
    .X(_14534_));
 sky130_fd_sc_hd__mux2_1 _18562_ (.A0(_14486_),
    .A1(\cpuregs[8][7] ),
    .S(_14534_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _18563_ (.A0(_14488_),
    .A1(\cpuregs[8][6] ),
    .S(_14534_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _18564_ (.A0(_14489_),
    .A1(\cpuregs[8][5] ),
    .S(_14534_),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_1 _18565_ (.A0(_14490_),
    .A1(\cpuregs[8][4] ),
    .S(_14534_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _18566_ (.A0(_14491_),
    .A1(\cpuregs[8][3] ),
    .S(_14534_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _18567_ (.A0(_14492_),
    .A1(\cpuregs[8][2] ),
    .S(_14534_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _18568_ (.A0(_14493_),
    .A1(\cpuregs[8][1] ),
    .S(_14529_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _18569_ (.A0(_14494_),
    .A1(\cpuregs[8][0] ),
    .S(_14529_),
    .X(_02771_));
 sky130_vsdinv _18570_ (.A(\reg_next_pc[0] ),
    .Y(_14535_));
 sky130_fd_sc_hd__buf_2 _18571_ (.A(latched_branch),
    .X(_14536_));
 sky130_fd_sc_hd__clkbuf_4 _18572_ (.A(latched_branch),
    .X(_14537_));
 sky130_fd_sc_hd__nor2_8 _18573_ (.A(_14537_),
    .B(_12863_),
    .Y(_00292_));
 sky130_fd_sc_hd__a211oi_4 _18574_ (.A1(_13736_),
    .A2(_14536_),
    .B1(_13101_),
    .C1(_00292_),
    .Y(_14538_));
 sky130_fd_sc_hd__nor3_1 _18575_ (.A(_13717_),
    .B(_14535_),
    .C(_14538_),
    .Y(_02770_));
 sky130_fd_sc_hd__clkbuf_2 _18576_ (.A(_12655_),
    .X(_14539_));
 sky130_fd_sc_hd__and2_1 _18577_ (.A(_14539_),
    .B(_00008_),
    .X(_02769_));
 sky130_fd_sc_hd__and2_1 _18578_ (.A(_14539_),
    .B(_15245_),
    .X(_02768_));
 sky130_fd_sc_hd__and2_1 _18579_ (.A(_14539_),
    .B(_00031_),
    .X(_02767_));
 sky130_fd_sc_hd__and2_1 _18580_ (.A(_14539_),
    .B(_00032_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_1 _18581_ (.A(_14539_),
    .B(_00033_),
    .X(_02765_));
 sky130_fd_sc_hd__and2_1 _18582_ (.A(_14539_),
    .B(_00034_),
    .X(_02764_));
 sky130_fd_sc_hd__buf_2 _18583_ (.A(_12655_),
    .X(_14540_));
 sky130_fd_sc_hd__and2_1 _18584_ (.A(_14540_),
    .B(_00035_),
    .X(_02763_));
 sky130_fd_sc_hd__and2_1 _18585_ (.A(_14540_),
    .B(_00036_),
    .X(_02762_));
 sky130_fd_sc_hd__and2_1 _18586_ (.A(_14540_),
    .B(_00037_),
    .X(_02761_));
 sky130_fd_sc_hd__and2_1 _18587_ (.A(_14540_),
    .B(_00009_),
    .X(_02760_));
 sky130_fd_sc_hd__and2_1 _18588_ (.A(_14540_),
    .B(_00010_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_1 _18589_ (.A(_14540_),
    .B(_00011_),
    .X(_02758_));
 sky130_fd_sc_hd__buf_2 _18590_ (.A(_12655_),
    .X(_14541_));
 sky130_fd_sc_hd__and2_1 _18591_ (.A(_14541_),
    .B(_00012_),
    .X(_02757_));
 sky130_fd_sc_hd__and2_1 _18592_ (.A(_14541_),
    .B(_00013_),
    .X(_02756_));
 sky130_fd_sc_hd__and2_1 _18593_ (.A(_14541_),
    .B(_00014_),
    .X(_02755_));
 sky130_fd_sc_hd__and2_1 _18594_ (.A(_14541_),
    .B(_00015_),
    .X(_02754_));
 sky130_fd_sc_hd__and2_1 _18595_ (.A(_14541_),
    .B(_00016_),
    .X(_02753_));
 sky130_fd_sc_hd__and2_1 _18596_ (.A(_14541_),
    .B(_00017_),
    .X(_02752_));
 sky130_fd_sc_hd__buf_2 _18597_ (.A(_12655_),
    .X(_14542_));
 sky130_fd_sc_hd__and2_1 _18598_ (.A(_14542_),
    .B(_00018_),
    .X(_02751_));
 sky130_fd_sc_hd__and2_1 _18599_ (.A(_14542_),
    .B(_00019_),
    .X(_02750_));
 sky130_fd_sc_hd__and2_1 _18600_ (.A(_14542_),
    .B(_00020_),
    .X(_02749_));
 sky130_fd_sc_hd__and2_1 _18601_ (.A(_14542_),
    .B(_00021_),
    .X(_02748_));
 sky130_fd_sc_hd__and2_1 _18602_ (.A(_14542_),
    .B(_00022_),
    .X(_02747_));
 sky130_fd_sc_hd__and2_1 _18603_ (.A(_14542_),
    .B(_00023_),
    .X(_02746_));
 sky130_fd_sc_hd__buf_2 _18604_ (.A(_12655_),
    .X(_14543_));
 sky130_fd_sc_hd__and2_1 _18605_ (.A(_14543_),
    .B(_00024_),
    .X(_02745_));
 sky130_fd_sc_hd__and2_1 _18606_ (.A(_14543_),
    .B(_00025_),
    .X(_02744_));
 sky130_fd_sc_hd__and2_1 _18607_ (.A(_14543_),
    .B(_00026_),
    .X(_02743_));
 sky130_fd_sc_hd__and2_1 _18608_ (.A(_14543_),
    .B(_00027_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_1 _18609_ (.A(_14543_),
    .B(_00028_),
    .X(_02741_));
 sky130_fd_sc_hd__and2_1 _18610_ (.A(_14543_),
    .B(_00029_),
    .X(_02740_));
 sky130_fd_sc_hd__and2_1 _18611_ (.A(_12650_),
    .B(_00030_),
    .X(_02739_));
 sky130_fd_sc_hd__nand2_1 _18612_ (.A(\decoded_imm_uj[1] ),
    .B(_12899_),
    .Y(_14544_));
 sky130_fd_sc_hd__o21ai_1 _18613_ (.A1(_12979_),
    .A2(_14111_),
    .B1(\mem_rdata_q[8] ),
    .Y(_14545_));
 sky130_fd_sc_hd__o211ai_1 _18614_ (.A1(_14172_),
    .A2(_14134_),
    .B1(_14544_),
    .C1(_14545_),
    .Y(_14546_));
 sky130_fd_sc_hd__mux2_1 _18615_ (.A0(_14546_),
    .A1(\decoded_imm[1] ),
    .S(_14136_),
    .X(_02738_));
 sky130_fd_sc_hd__nand2_1 _18616_ (.A(\decoded_imm_uj[2] ),
    .B(_12899_),
    .Y(_14547_));
 sky130_fd_sc_hd__o21ai_1 _18617_ (.A1(_12979_),
    .A2(_14111_),
    .B1(\mem_rdata_q[9] ),
    .Y(_14548_));
 sky130_fd_sc_hd__o211ai_1 _18618_ (.A1(_14165_),
    .A2(_14134_),
    .B1(_14547_),
    .C1(_14548_),
    .Y(_14549_));
 sky130_fd_sc_hd__mux2_1 _18619_ (.A0(_14549_),
    .A1(\decoded_imm[2] ),
    .S(_14136_),
    .X(_02737_));
 sky130_fd_sc_hd__nand2_1 _18620_ (.A(\decoded_imm_uj[3] ),
    .B(_12899_),
    .Y(_14550_));
 sky130_fd_sc_hd__o21ai_1 _18621_ (.A1(_12979_),
    .A2(_14111_),
    .B1(\mem_rdata_q[10] ),
    .Y(_14551_));
 sky130_fd_sc_hd__o211ai_1 _18622_ (.A1(_14164_),
    .A2(_14134_),
    .B1(_14550_),
    .C1(_14551_),
    .Y(_14552_));
 sky130_fd_sc_hd__mux2_1 _18623_ (.A0(_14552_),
    .A1(\decoded_imm[3] ),
    .S(_14136_),
    .X(_02736_));
 sky130_vsdinv _18624_ (.A(\decoded_imm[4] ),
    .Y(_14553_));
 sky130_fd_sc_hd__inv_2 _18625_ (.A(\decoded_imm_uj[4] ),
    .Y(_00367_));
 sky130_vsdinv _18626_ (.A(\mem_rdata_q[24] ),
    .Y(_14554_));
 sky130_fd_sc_hd__o21ai_1 _18627_ (.A1(_12978_),
    .A2(_14111_),
    .B1(\mem_rdata_q[11] ),
    .Y(_14555_));
 sky130_fd_sc_hd__o221a_1 _18628_ (.A1(_00367_),
    .A2(_12821_),
    .B1(_14554_),
    .B2(_14133_),
    .C1(_14555_),
    .X(_14556_));
 sky130_fd_sc_hd__or2b_1 _18629_ (.A(_14556_),
    .B_N(_13070_),
    .X(_14557_));
 sky130_fd_sc_hd__o21ai_1 _18630_ (.A1(_14553_),
    .A2(_14113_),
    .B1(_14557_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand3_4 _18631_ (.A(_14133_),
    .B(_13571_),
    .C(_12884_),
    .Y(_14558_));
 sky130_fd_sc_hd__clkbuf_2 _18632_ (.A(_14558_),
    .X(_14559_));
 sky130_vsdinv _18633_ (.A(\decoded_imm_uj[5] ),
    .Y(_14560_));
 sky130_fd_sc_hd__o2bb2ai_1 _18634_ (.A1_N(_14154_),
    .A2_N(_14559_),
    .B1(_14560_),
    .B2(_00323_),
    .Y(_14561_));
 sky130_fd_sc_hd__mux2_1 _18635_ (.A0(_14561_),
    .A1(\decoded_imm[5] ),
    .S(_14136_),
    .X(_02734_));
 sky130_fd_sc_hd__a22o_1 _18636_ (.A1(\decoded_imm_uj[6] ),
    .A2(_12900_),
    .B1(_14559_),
    .B2(\mem_rdata_q[26] ),
    .X(_14562_));
 sky130_fd_sc_hd__clkbuf_4 _18637_ (.A(\decoded_imm[6] ),
    .X(_14563_));
 sky130_fd_sc_hd__mux2_1 _18638_ (.A0(_14562_),
    .A1(_14563_),
    .S(_14136_),
    .X(_02733_));
 sky130_vsdinv _18639_ (.A(\decoded_imm_uj[7] ),
    .Y(_14564_));
 sky130_fd_sc_hd__o2bb2ai_1 _18640_ (.A1_N(_14141_),
    .A2_N(_14559_),
    .B1(_14564_),
    .B2(_00323_),
    .Y(_14565_));
 sky130_fd_sc_hd__clkbuf_2 _18641_ (.A(\decoded_imm[7] ),
    .X(_14566_));
 sky130_fd_sc_hd__buf_2 _18642_ (.A(_13004_),
    .X(_14567_));
 sky130_fd_sc_hd__mux2_1 _18643_ (.A0(_14565_),
    .A1(_14566_),
    .S(_14567_),
    .X(_02732_));
 sky130_fd_sc_hd__a22o_1 _18644_ (.A1(\decoded_imm_uj[8] ),
    .A2(_12900_),
    .B1(_14559_),
    .B2(\mem_rdata_q[28] ),
    .X(_14568_));
 sky130_fd_sc_hd__clkbuf_4 _18645_ (.A(\decoded_imm[8] ),
    .X(_14569_));
 sky130_fd_sc_hd__mux2_1 _18646_ (.A0(_14568_),
    .A1(_14569_),
    .S(_14567_),
    .X(_02731_));
 sky130_fd_sc_hd__a22o_1 _18647_ (.A1(\decoded_imm_uj[9] ),
    .A2(_12900_),
    .B1(_14559_),
    .B2(_13014_),
    .X(_14570_));
 sky130_fd_sc_hd__buf_2 _18648_ (.A(\decoded_imm[9] ),
    .X(_14571_));
 sky130_fd_sc_hd__mux2_1 _18649_ (.A0(_14570_),
    .A1(_14571_),
    .S(_14567_),
    .X(_02730_));
 sky130_fd_sc_hd__clkbuf_2 _18650_ (.A(_14558_),
    .X(_14572_));
 sky130_fd_sc_hd__a22o_1 _18651_ (.A1(\decoded_imm_uj[10] ),
    .A2(_12900_),
    .B1(_14572_),
    .B2(\mem_rdata_q[30] ),
    .X(_14573_));
 sky130_fd_sc_hd__mux2_1 _18652_ (.A0(_14573_),
    .A1(\decoded_imm[10] ),
    .S(_14567_),
    .X(_02729_));
 sky130_vsdinv _18653_ (.A(\decoded_imm[11] ),
    .Y(_14574_));
 sky130_fd_sc_hd__nand2_1 _18654_ (.A(_14134_),
    .B(_12884_),
    .Y(_14575_));
 sky130_fd_sc_hd__and2_1 _18655_ (.A(_12978_),
    .B(\mem_rdata_q[7] ),
    .X(_14576_));
 sky130_fd_sc_hd__a221oi_2 _18656_ (.A1(\decoded_imm_uj[11] ),
    .A2(_12899_),
    .B1(_14575_),
    .B2(_14206_),
    .C1(_14576_),
    .Y(_14577_));
 sky130_fd_sc_hd__or2b_1 _18657_ (.A(_14577_),
    .B_N(_13070_),
    .X(_14578_));
 sky130_fd_sc_hd__o21ai_1 _18658_ (.A1(_14574_),
    .A2(_14113_),
    .B1(_14578_),
    .Y(_02728_));
 sky130_vsdinv _18659_ (.A(_12820_),
    .Y(_14579_));
 sky130_fd_sc_hd__clkbuf_2 _18660_ (.A(_14579_),
    .X(_14580_));
 sky130_fd_sc_hd__and2_1 _18661_ (.A(\decoded_imm_uj[12] ),
    .B(_12899_),
    .X(_14581_));
 sky130_fd_sc_hd__a221o_1 _18662_ (.A1(_12994_),
    .A2(_14580_),
    .B1(_14572_),
    .B2(_14207_),
    .C1(_14581_),
    .X(_14582_));
 sky130_fd_sc_hd__mux2_1 _18663_ (.A0(_14582_),
    .A1(\decoded_imm[12] ),
    .S(_14567_),
    .X(_02727_));
 sky130_fd_sc_hd__buf_1 _18664_ (.A(instr_jal),
    .X(_14583_));
 sky130_fd_sc_hd__and2_1 _18665_ (.A(\decoded_imm_uj[13] ),
    .B(_14583_),
    .X(_14584_));
 sky130_fd_sc_hd__a221o_1 _18666_ (.A1(_12992_),
    .A2(_14580_),
    .B1(_14572_),
    .B2(_14207_),
    .C1(_14584_),
    .X(_14585_));
 sky130_fd_sc_hd__mux2_1 _18667_ (.A0(_14585_),
    .A1(\decoded_imm[13] ),
    .S(_14567_),
    .X(_02726_));
 sky130_vsdinv _18668_ (.A(\decoded_imm_uj[14] ),
    .Y(_14586_));
 sky130_fd_sc_hd__nand2_1 _18669_ (.A(_14572_),
    .B(_14207_),
    .Y(_14587_));
 sky130_fd_sc_hd__o221ai_2 _18670_ (.A1(_14586_),
    .A2(_12821_),
    .B1(_00334_),
    .B2(_12820_),
    .C1(_14587_),
    .Y(_14588_));
 sky130_fd_sc_hd__buf_2 _18671_ (.A(_13004_),
    .X(_14589_));
 sky130_fd_sc_hd__mux2_1 _18672_ (.A0(_14588_),
    .A1(\decoded_imm[14] ),
    .S(_14589_),
    .X(_02725_));
 sky130_fd_sc_hd__and2_1 _18673_ (.A(\decoded_imm_uj[15] ),
    .B(_14583_),
    .X(_14590_));
 sky130_fd_sc_hd__a221o_1 _18674_ (.A1(\mem_rdata_q[15] ),
    .A2(_14580_),
    .B1(_14572_),
    .B2(_14207_),
    .C1(_14590_),
    .X(_14591_));
 sky130_fd_sc_hd__mux2_1 _18675_ (.A0(_14591_),
    .A1(\decoded_imm[15] ),
    .S(_14589_),
    .X(_02724_));
 sky130_fd_sc_hd__and2_1 _18676_ (.A(\decoded_imm_uj[16] ),
    .B(_14583_),
    .X(_14592_));
 sky130_fd_sc_hd__a221o_1 _18677_ (.A1(\mem_rdata_q[16] ),
    .A2(_14580_),
    .B1(_14572_),
    .B2(_14206_),
    .C1(_14592_),
    .X(_14593_));
 sky130_fd_sc_hd__buf_2 _18678_ (.A(\decoded_imm[16] ),
    .X(_14594_));
 sky130_fd_sc_hd__mux2_1 _18679_ (.A0(_14593_),
    .A1(_14594_),
    .S(_14589_),
    .X(_02723_));
 sky130_fd_sc_hd__and2_1 _18680_ (.A(\decoded_imm_uj[17] ),
    .B(_14583_),
    .X(_14595_));
 sky130_fd_sc_hd__a221o_1 _18681_ (.A1(\mem_rdata_q[17] ),
    .A2(_14580_),
    .B1(_14558_),
    .B2(_14206_),
    .C1(_14595_),
    .X(_14596_));
 sky130_fd_sc_hd__clkbuf_4 _18682_ (.A(\decoded_imm[17] ),
    .X(_14597_));
 sky130_fd_sc_hd__mux2_1 _18683_ (.A0(_14596_),
    .A1(_14597_),
    .S(_14589_),
    .X(_02722_));
 sky130_fd_sc_hd__and2_1 _18684_ (.A(\decoded_imm_uj[18] ),
    .B(_14583_),
    .X(_14598_));
 sky130_fd_sc_hd__a221o_1 _18685_ (.A1(\mem_rdata_q[18] ),
    .A2(_14580_),
    .B1(_14558_),
    .B2(_14206_),
    .C1(_14598_),
    .X(_14599_));
 sky130_fd_sc_hd__clkbuf_4 _18686_ (.A(\decoded_imm[18] ),
    .X(_14600_));
 sky130_fd_sc_hd__mux2_1 _18687_ (.A0(_14599_),
    .A1(_14600_),
    .S(_14589_),
    .X(_02721_));
 sky130_fd_sc_hd__and2_1 _18688_ (.A(\decoded_imm_uj[19] ),
    .B(_14583_),
    .X(_14601_));
 sky130_fd_sc_hd__a221o_1 _18689_ (.A1(\mem_rdata_q[19] ),
    .A2(_14579_),
    .B1(_14558_),
    .B2(_14206_),
    .C1(_14601_),
    .X(_14602_));
 sky130_fd_sc_hd__mux2_1 _18690_ (.A0(_14602_),
    .A1(\decoded_imm[19] ),
    .S(_14589_),
    .X(_02720_));
 sky130_fd_sc_hd__nor2_4 _18691_ (.A(_14177_),
    .B(_14134_),
    .Y(_14603_));
 sky130_fd_sc_hd__clkbuf_2 _18692_ (.A(_14603_),
    .X(_14604_));
 sky130_fd_sc_hd__buf_2 _18693_ (.A(_14579_),
    .X(_14605_));
 sky130_fd_sc_hd__clkbuf_2 _18694_ (.A(_13004_),
    .X(_14606_));
 sky130_fd_sc_hd__nor2_1 _18695_ (.A(_12978_),
    .B(is_sb_sh_sw),
    .Y(_14607_));
 sky130_fd_sc_hd__o2bb2ai_2 _18696_ (.A1_N(_14126_),
    .A2_N(instr_jal),
    .B1(_14177_),
    .B2(_14607_),
    .Y(_14608_));
 sky130_fd_sc_hd__buf_2 _18697_ (.A(_14608_),
    .X(_14609_));
 sky130_fd_sc_hd__a211o_1 _18698_ (.A1(\mem_rdata_q[20] ),
    .A2(_14605_),
    .B1(_14606_),
    .C1(_14609_),
    .X(_14610_));
 sky130_fd_sc_hd__o22a_1 _18699_ (.A1(\decoded_imm[20] ),
    .A2(_13572_),
    .B1(_14604_),
    .B2(_14610_),
    .X(_02719_));
 sky130_fd_sc_hd__a211o_1 _18700_ (.A1(\mem_rdata_q[21] ),
    .A2(_14605_),
    .B1(_14606_),
    .C1(_14609_),
    .X(_14611_));
 sky130_fd_sc_hd__o22a_1 _18701_ (.A1(\decoded_imm[21] ),
    .A2(_13572_),
    .B1(_14604_),
    .B2(_14611_),
    .X(_02718_));
 sky130_fd_sc_hd__a211o_1 _18702_ (.A1(\mem_rdata_q[22] ),
    .A2(_14605_),
    .B1(_14606_),
    .C1(_14609_),
    .X(_14612_));
 sky130_fd_sc_hd__o22a_1 _18703_ (.A1(\decoded_imm[22] ),
    .A2(_13572_),
    .B1(_14604_),
    .B2(_14612_),
    .X(_02717_));
 sky130_fd_sc_hd__clkbuf_2 _18704_ (.A(_14157_),
    .X(_14613_));
 sky130_fd_sc_hd__a211o_1 _18705_ (.A1(\mem_rdata_q[23] ),
    .A2(_14605_),
    .B1(_14606_),
    .C1(_14609_),
    .X(_14614_));
 sky130_fd_sc_hd__o22a_1 _18706_ (.A1(\decoded_imm[23] ),
    .A2(_14613_),
    .B1(_14604_),
    .B2(_14614_),
    .X(_02716_));
 sky130_fd_sc_hd__buf_4 _18707_ (.A(\decoded_imm[24] ),
    .X(_14615_));
 sky130_fd_sc_hd__clkbuf_2 _18708_ (.A(_14579_),
    .X(_14616_));
 sky130_fd_sc_hd__a211o_1 _18709_ (.A1(\mem_rdata_q[24] ),
    .A2(_14616_),
    .B1(_14606_),
    .C1(_14608_),
    .X(_14617_));
 sky130_fd_sc_hd__o22a_1 _18710_ (.A1(_14615_),
    .A2(_14613_),
    .B1(_14604_),
    .B2(_14617_),
    .X(_02715_));
 sky130_fd_sc_hd__clkbuf_4 _18711_ (.A(\decoded_imm[25] ),
    .X(_14618_));
 sky130_fd_sc_hd__a211o_1 _18712_ (.A1(_14154_),
    .A2(_14616_),
    .B1(_14606_),
    .C1(_14608_),
    .X(_14619_));
 sky130_fd_sc_hd__o22a_1 _18713_ (.A1(_14618_),
    .A2(_14613_),
    .B1(_14604_),
    .B2(_14619_),
    .X(_02714_));
 sky130_fd_sc_hd__buf_2 _18714_ (.A(\decoded_imm[26] ),
    .X(_14620_));
 sky130_vsdinv _18715_ (.A(_14620_),
    .Y(_14621_));
 sky130_fd_sc_hd__a2111oi_2 _18716_ (.A1(\mem_rdata_q[26] ),
    .A2(_14605_),
    .B1(_13056_),
    .C1(_14609_),
    .D1(_14603_),
    .Y(_14622_));
 sky130_fd_sc_hd__a21oi_1 _18717_ (.A1(_14621_),
    .A2(_14156_),
    .B1(_14622_),
    .Y(_02713_));
 sky130_fd_sc_hd__buf_2 _18718_ (.A(\decoded_imm[27] ),
    .X(_14623_));
 sky130_fd_sc_hd__a211o_1 _18719_ (.A1(_14141_),
    .A2(_14616_),
    .B1(_13059_),
    .C1(_14608_),
    .X(_14624_));
 sky130_fd_sc_hd__o22a_1 _18720_ (.A1(_14623_),
    .A2(_14613_),
    .B1(_14603_),
    .B2(_14624_),
    .X(_02712_));
 sky130_fd_sc_hd__buf_2 _18721_ (.A(\decoded_imm[28] ),
    .X(_14625_));
 sky130_fd_sc_hd__a211o_1 _18722_ (.A1(\mem_rdata_q[28] ),
    .A2(_14616_),
    .B1(_13059_),
    .C1(_14608_),
    .X(_14626_));
 sky130_fd_sc_hd__o22a_1 _18723_ (.A1(_14625_),
    .A2(_14613_),
    .B1(_14603_),
    .B2(_14626_),
    .X(_02711_));
 sky130_vsdinv _18724_ (.A(\decoded_imm[29] ),
    .Y(_14627_));
 sky130_fd_sc_hd__a2111oi_2 _18725_ (.A1(_13014_),
    .A2(_14605_),
    .B1(_13056_),
    .C1(_14609_),
    .D1(_14603_),
    .Y(_14628_));
 sky130_fd_sc_hd__a21oi_1 _18726_ (.A1(_14627_),
    .A2(_14156_),
    .B1(_14628_),
    .Y(_02710_));
 sky130_fd_sc_hd__a211o_1 _18727_ (.A1(\mem_rdata_q[30] ),
    .A2(_14616_),
    .B1(_13059_),
    .C1(_14608_),
    .X(_14629_));
 sky130_fd_sc_hd__o22a_1 _18728_ (.A1(\decoded_imm[30] ),
    .A2(_14613_),
    .B1(_14603_),
    .B2(_14629_),
    .X(_02709_));
 sky130_fd_sc_hd__clkinv_8 _18729_ (.A(\decoded_imm_uj[20] ),
    .Y(_14630_));
 sky130_fd_sc_hd__nor2_1 _18730_ (.A(_14616_),
    .B(_14559_),
    .Y(_14631_));
 sky130_fd_sc_hd__o22ai_2 _18731_ (.A1(_14630_),
    .A2(_00323_),
    .B1(_14177_),
    .B2(_14631_),
    .Y(_14632_));
 sky130_fd_sc_hd__mux2_1 _18732_ (.A0(_14632_),
    .A1(\decoded_imm[31] ),
    .S(_13056_),
    .X(_02708_));
 sky130_fd_sc_hd__o311a_4 _18733_ (.A1(_12978_),
    .A2(_12846_),
    .A3(_12811_),
    .B1(_12852_),
    .C1(_13873_),
    .X(_14633_));
 sky130_fd_sc_hd__nor2_8 _18734_ (.A(_12845_),
    .B(_12915_),
    .Y(_14634_));
 sky130_fd_sc_hd__nand3_4 _18735_ (.A(_14633_),
    .B(_15205_),
    .C(_14634_),
    .Y(_14635_));
 sky130_fd_sc_hd__o21ai_1 _18736_ (.A1(_13785_),
    .A2(_14633_),
    .B1(_14635_),
    .Y(_02707_));
 sky130_vsdinv _18737_ (.A(_14634_),
    .Y(_02542_));
 sky130_vsdinv _18738_ (.A(_14633_),
    .Y(_14636_));
 sky130_fd_sc_hd__and4_4 _18739_ (.A(_12771_),
    .B(_12873_),
    .C(_14633_),
    .D(_14634_),
    .X(_14637_));
 sky130_fd_sc_hd__a22o_1 _18740_ (.A1(\latched_rd[1] ),
    .A2(_14636_),
    .B1(_14637_),
    .B2(\decoded_rd[1] ),
    .X(_02706_));
 sky130_fd_sc_hd__a22o_1 _18741_ (.A1(_13745_),
    .A2(_14636_),
    .B1(_14637_),
    .B2(\decoded_rd[2] ),
    .X(_02705_));
 sky130_fd_sc_hd__a22o_1 _18742_ (.A1(_13744_),
    .A2(_14636_),
    .B1(_14637_),
    .B2(\decoded_rd[3] ),
    .X(_02704_));
 sky130_vsdinv _18743_ (.A(_12842_),
    .Y(_14638_));
 sky130_fd_sc_hd__nor3_1 _18744_ (.A(_14111_),
    .B(_14638_),
    .C(_00310_),
    .Y(_14639_));
 sky130_vsdinv _18745_ (.A(_14639_),
    .Y(_14640_));
 sky130_fd_sc_hd__o31ai_4 _18746_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(is_slli_srli_srai),
    .A3(is_lui_auipc_jal),
    .B1(_12916_),
    .Y(_14641_));
 sky130_fd_sc_hd__a21oi_1 _18747_ (.A1(_14640_),
    .A2(_14641_),
    .B1(_13796_),
    .Y(_02703_));
 sky130_fd_sc_hd__buf_2 _18748_ (.A(_13832_),
    .X(_14642_));
 sky130_fd_sc_hd__nor2b_1 _18749_ (.A(_14642_),
    .B_N(_02558_),
    .Y(_02702_));
 sky130_fd_sc_hd__nor2b_1 _18750_ (.A(_14642_),
    .B_N(_02557_),
    .Y(_02701_));
 sky130_fd_sc_hd__nor2b_1 _18751_ (.A(_14642_),
    .B_N(_02556_),
    .Y(_02700_));
 sky130_fd_sc_hd__nor2b_1 _18752_ (.A(_14642_),
    .B_N(_02555_),
    .Y(_02699_));
 sky130_fd_sc_hd__nor2b_1 _18753_ (.A(_14642_),
    .B_N(_02554_),
    .Y(_02698_));
 sky130_fd_sc_hd__nor2b_1 _18754_ (.A(_14642_),
    .B_N(_02553_),
    .Y(_02697_));
 sky130_fd_sc_hd__buf_2 _18755_ (.A(_13831_),
    .X(_14643_));
 sky130_fd_sc_hd__nor2b_1 _18756_ (.A(_14643_),
    .B_N(_02552_),
    .Y(_02696_));
 sky130_fd_sc_hd__nor2b_1 _18757_ (.A(_14643_),
    .B_N(_02551_),
    .Y(_02695_));
 sky130_fd_sc_hd__buf_2 _18758_ (.A(_13834_),
    .X(_14644_));
 sky130_fd_sc_hd__nor2b_1 _18759_ (.A(_14644_),
    .B_N(_00122_),
    .Y(_02550_));
 sky130_fd_sc_hd__clkbuf_4 _18760_ (.A(_13834_),
    .X(_14645_));
 sky130_fd_sc_hd__nor3b_1 _18761_ (.A(_14643_),
    .B(_14645_),
    .C_N(_00122_),
    .Y(_02694_));
 sky130_fd_sc_hd__nor2b_1 _18762_ (.A(_14644_),
    .B_N(_00116_),
    .Y(_02549_));
 sky130_fd_sc_hd__nor3b_1 _18763_ (.A(_14643_),
    .B(_14645_),
    .C_N(_00116_),
    .Y(_02693_));
 sky130_fd_sc_hd__nor2b_1 _18764_ (.A(_14644_),
    .B_N(_00110_),
    .Y(_02548_));
 sky130_fd_sc_hd__nor3b_1 _18765_ (.A(_14643_),
    .B(_14645_),
    .C_N(_00110_),
    .Y(_02692_));
 sky130_fd_sc_hd__nor2b_1 _18766_ (.A(_14644_),
    .B_N(_00104_),
    .Y(_02547_));
 sky130_fd_sc_hd__nor3b_1 _18767_ (.A(_13832_),
    .B(_14645_),
    .C_N(_00104_),
    .Y(_02691_));
 sky130_fd_sc_hd__clkbuf_4 _18768_ (.A(_13836_),
    .X(_14646_));
 sky130_fd_sc_hd__nor3b_1 _18769_ (.A(_14644_),
    .B(_14646_),
    .C_N(_00094_),
    .Y(_02546_));
 sky130_vsdinv _18770_ (.A(_13831_),
    .Y(_14647_));
 sky130_fd_sc_hd__clkbuf_2 _18771_ (.A(_14647_),
    .X(_02327_));
 sky130_vsdinv _18772_ (.A(net225),
    .Y(_14648_));
 sky130_fd_sc_hd__buf_1 _18773_ (.A(_14648_),
    .X(_02324_));
 sky130_vsdinv _18774_ (.A(net222),
    .Y(_14649_));
 sky130_fd_sc_hd__buf_1 _18775_ (.A(_14649_),
    .X(_02321_));
 sky130_fd_sc_hd__and4_1 _18776_ (.A(_02327_),
    .B(_02324_),
    .C(_02321_),
    .D(_00094_),
    .X(_02690_));
 sky130_fd_sc_hd__nor3b_2 _18777_ (.A(_14645_),
    .B(_14646_),
    .C_N(_00084_),
    .Y(_02545_));
 sky130_fd_sc_hd__and4_1 _18778_ (.A(_02327_),
    .B(_02324_),
    .C(_14649_),
    .D(_00084_),
    .X(_02689_));
 sky130_fd_sc_hd__inv_2 _18779_ (.A(net492),
    .Y(_02318_));
 sky130_fd_sc_hd__and4_1 _18780_ (.A(_02324_),
    .B(_02321_),
    .C(_02318_),
    .D(_00066_),
    .X(_02544_));
 sky130_fd_sc_hd__nor2b_2 _18781_ (.A(_13837_),
    .B_N(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__and4_1 _18782_ (.A(_00067_),
    .B(_02327_),
    .C(_02324_),
    .D(_02321_),
    .X(_02688_));
 sky130_fd_sc_hd__nor2b_2 _18783_ (.A(_13839_),
    .B_N(net306),
    .Y(_00048_));
 sky130_fd_sc_hd__and4_1 _18784_ (.A(_00048_),
    .B(_02324_),
    .C(_14649_),
    .D(_02318_),
    .X(_02543_));
 sky130_fd_sc_hd__nor3b_4 _18785_ (.A(net492),
    .B(_13839_),
    .C_N(_14266_),
    .Y(_00049_));
 sky130_fd_sc_hd__and4_1 _18786_ (.A(_00049_),
    .B(_02327_),
    .C(_14648_),
    .D(_02321_),
    .X(_02687_));
 sky130_fd_sc_hd__o211a_1 _18787_ (.A1(\reg_pc[1] ),
    .A2(\reg_next_pc[0] ),
    .B1(net101),
    .C1(mem_do_rinst),
    .X(_14650_));
 sky130_fd_sc_hd__clkbuf_2 _18788_ (.A(_14650_),
    .X(_00307_));
 sky130_fd_sc_hd__clkbuf_2 _18789_ (.A(irq_active),
    .X(_14651_));
 sky130_fd_sc_hd__nor3_1 _18790_ (.A(_14651_),
    .B(_12971_),
    .C(_13537_),
    .Y(_00312_));
 sky130_fd_sc_hd__o21a_1 _18791_ (.A1(mem_do_wdata),
    .A2(_12645_),
    .B1(net101),
    .X(_00303_));
 sky130_fd_sc_hd__nand3b_4 _18792_ (.A_N(_12997_),
    .B(_12774_),
    .C(_12674_),
    .Y(_14652_));
 sky130_fd_sc_hd__nor3_1 _18793_ (.A(irq_active),
    .B(_13540_),
    .C(\pcpi_mul.active[1] ),
    .Y(_14653_));
 sky130_fd_sc_hd__o21a_1 _18794_ (.A1(instr_ecall_ebreak),
    .A2(pcpi_timeout),
    .B1(_14653_),
    .X(_14654_));
 sky130_fd_sc_hd__nand3_4 _18795_ (.A(_00310_),
    .B(_12842_),
    .C(_14654_),
    .Y(_14655_));
 sky130_fd_sc_hd__o32ai_4 _18796_ (.A1(_12848_),
    .A2(_00309_),
    .A3(_14652_),
    .B1(_12643_),
    .B2(_14655_),
    .Y(_14656_));
 sky130_vsdinv _18797_ (.A(_00307_),
    .Y(_14657_));
 sky130_fd_sc_hd__clkbuf_4 _18798_ (.A(\mem_wordsize[2] ),
    .X(_14658_));
 sky130_fd_sc_hd__nor2_4 _18799_ (.A(irq_active),
    .B(\irq_mask[2] ),
    .Y(_14659_));
 sky130_fd_sc_hd__buf_2 _18800_ (.A(_14659_),
    .X(_14660_));
 sky130_fd_sc_hd__and4_1 _18801_ (.A(_14657_),
    .B(_14267_),
    .C(_14658_),
    .D(_14660_),
    .X(_14661_));
 sky130_fd_sc_hd__nor2_4 _18802_ (.A(_13565_),
    .B(_13566_),
    .Y(_14662_));
 sky130_fd_sc_hd__and3_1 _18803_ (.A(_14662_),
    .B(_12875_),
    .C(_14661_),
    .X(_14663_));
 sky130_fd_sc_hd__and2_1 _18804_ (.A(_14266_),
    .B(\mem_wordsize[2] ),
    .X(_14664_));
 sky130_fd_sc_hd__buf_2 _18805_ (.A(_14664_),
    .X(_00306_));
 sky130_fd_sc_hd__o21a_2 _18806_ (.A1(_14263_),
    .A2(_14266_),
    .B1(\mem_wordsize[0] ),
    .X(_00305_));
 sky130_fd_sc_hd__nor2_2 _18807_ (.A(_00306_),
    .B(_00305_),
    .Y(_14665_));
 sky130_fd_sc_hd__o211a_1 _18808_ (.A1(_14660_),
    .A2(_14665_),
    .B1(_14657_),
    .C1(_03828_),
    .X(_14666_));
 sky130_fd_sc_hd__a211o_1 _18809_ (.A1(_14656_),
    .A2(_14661_),
    .B1(_14663_),
    .C1(_14666_),
    .X(_14667_));
 sky130_vsdinv _18810_ (.A(_00303_),
    .Y(_14668_));
 sky130_fd_sc_hd__o21a_2 _18811_ (.A1(_14668_),
    .A2(_14665_),
    .B1(_14657_),
    .X(_14669_));
 sky130_fd_sc_hd__o21a_1 _18812_ (.A1(_14660_),
    .A2(_14669_),
    .B1(\pcpi_mul.active[1] ),
    .X(_14670_));
 sky130_fd_sc_hd__o2111a_1 _18813_ (.A1(\reg_pc[1] ),
    .A2(\reg_next_pc[0] ),
    .B1(_12638_),
    .C1(mem_do_rinst),
    .D1(_14659_),
    .X(_14671_));
 sky130_fd_sc_hd__nor2_1 _18814_ (.A(_14671_),
    .B(_14669_),
    .Y(_14672_));
 sky130_fd_sc_hd__a211oi_4 _18815_ (.A1(_14267_),
    .A2(_14658_),
    .B1(_12641_),
    .C1(_12635_),
    .Y(_14673_));
 sky130_fd_sc_hd__o211a_1 _18816_ (.A1(_14263_),
    .A2(_14266_),
    .B1(\mem_wordsize[0] ),
    .C1(_14659_),
    .X(_14674_));
 sky130_fd_sc_hd__nand3b_1 _18817_ (.A_N(_00307_),
    .B(_14673_),
    .C(_14674_),
    .Y(_14675_));
 sky130_fd_sc_hd__a21boi_1 _18818_ (.A1(_14672_),
    .A2(_14675_),
    .B1_N(_14654_),
    .Y(_14676_));
 sky130_fd_sc_hd__o2111a_1 _18819_ (.A1(_14670_),
    .A2(_14676_),
    .B1(_12843_),
    .C1(_12887_),
    .D1(_12886_),
    .X(_14677_));
 sky130_vsdinv _18820_ (.A(_14659_),
    .Y(_14678_));
 sky130_fd_sc_hd__nand2_1 _18821_ (.A(_14650_),
    .B(_14678_),
    .Y(_14679_));
 sky130_fd_sc_hd__o211a_1 _18822_ (.A1(_00307_),
    .A2(_14668_),
    .B1(_14679_),
    .C1(_03828_),
    .X(_14680_));
 sky130_fd_sc_hd__nor3_4 _18823_ (.A(net494),
    .B(_12832_),
    .C(_12854_),
    .Y(_14681_));
 sky130_fd_sc_hd__o221ai_2 _18824_ (.A1(mem_do_wdata),
    .A2(_12645_),
    .B1(_00306_),
    .B2(_00305_),
    .C1(_14678_),
    .Y(_14682_));
 sky130_fd_sc_hd__and3_1 _18825_ (.A(_14682_),
    .B(_12638_),
    .C(_14679_),
    .X(_14683_));
 sky130_vsdinv _18826_ (.A(_14683_),
    .Y(_14684_));
 sky130_fd_sc_hd__nand3b_1 _18827_ (.A_N(_12639_),
    .B(\cpu_state[4] ),
    .C(_12816_),
    .Y(_14685_));
 sky130_fd_sc_hd__o2bb2ai_1 _18828_ (.A1_N(_13875_),
    .A2_N(_14685_),
    .B1(_14660_),
    .B2(_14669_),
    .Y(_14686_));
 sky130_fd_sc_hd__o31ai_2 _18829_ (.A1(_12853_),
    .A2(_14681_),
    .A3(_14684_),
    .B1(_14686_),
    .Y(_14687_));
 sky130_fd_sc_hd__or4_4 _18830_ (.A(_12870_),
    .B(_00314_),
    .C(_14680_),
    .D(_14687_),
    .X(_14688_));
 sky130_vsdinv _18831_ (.A(_00305_),
    .Y(_14689_));
 sky130_fd_sc_hd__o2111ai_4 _18832_ (.A1(_14660_),
    .A2(_14689_),
    .B1(_14657_),
    .C1(_14673_),
    .D1(_14662_),
    .Y(_14690_));
 sky130_fd_sc_hd__o2111a_1 _18833_ (.A1(_12696_),
    .A2(_12697_),
    .B1(instr_jal),
    .C1(decoder_trigger),
    .D1(_12774_),
    .X(_02062_));
 sky130_fd_sc_hd__nand3_1 _18834_ (.A(_02062_),
    .B(_12674_),
    .C(_14674_),
    .Y(_14691_));
 sky130_fd_sc_hd__a2111o_1 _18835_ (.A1(instr_waitirq),
    .A2(do_waitirq),
    .B1(_12997_),
    .C1(_00305_),
    .D1(_13566_),
    .X(_14692_));
 sky130_fd_sc_hd__a21bo_1 _18836_ (.A1(_14691_),
    .A2(_14692_),
    .B1_N(_14673_),
    .X(_14693_));
 sky130_fd_sc_hd__a21oi_2 _18837_ (.A1(_14673_),
    .A2(_14674_),
    .B1(_14668_),
    .Y(_14694_));
 sky130_fd_sc_hd__a2111o_1 _18838_ (.A1(instr_waitirq),
    .A2(do_waitirq),
    .B1(_12997_),
    .C1(_14694_),
    .D1(_13566_),
    .X(_14695_));
 sky130_vsdinv _18839_ (.A(_12645_),
    .Y(_14696_));
 sky130_fd_sc_hd__a21o_1 _18840_ (.A1(_12771_),
    .A2(_12873_),
    .B1(_12641_),
    .X(_14697_));
 sky130_fd_sc_hd__a2111o_1 _18841_ (.A1(_00291_),
    .A2(_14696_),
    .B1(_14678_),
    .C1(_14665_),
    .D1(_14697_),
    .X(_14698_));
 sky130_fd_sc_hd__o21a_1 _18842_ (.A1(_12635_),
    .A2(_14665_),
    .B1(_12674_),
    .X(_14699_));
 sky130_fd_sc_hd__a22oi_1 _18843_ (.A1(_14662_),
    .A2(_14668_),
    .B1(_02062_),
    .B2(_14699_),
    .Y(_14700_));
 sky130_fd_sc_hd__a41o_1 _18844_ (.A1(_14693_),
    .A2(_14695_),
    .A3(_14698_),
    .A4(_14700_),
    .B1(_00307_),
    .X(_14701_));
 sky130_fd_sc_hd__a31oi_2 _18845_ (.A1(_14659_),
    .A2(_00303_),
    .A3(_00306_),
    .B1(_14671_),
    .Y(_14702_));
 sky130_fd_sc_hd__nand3b_1 _18846_ (.A_N(_14702_),
    .B(_02062_),
    .C(_12648_),
    .Y(_14703_));
 sky130_fd_sc_hd__o21a_1 _18847_ (.A1(_14697_),
    .A2(_14672_),
    .B1(_14703_),
    .X(_14704_));
 sky130_fd_sc_hd__a21bo_1 _18848_ (.A1(_14652_),
    .A2(_13565_),
    .B1_N(_14671_),
    .X(_14705_));
 sky130_fd_sc_hd__a41oi_1 _18849_ (.A1(_14690_),
    .A2(_14701_),
    .A3(_14704_),
    .A4(_14705_),
    .B1(_13101_),
    .Y(_14706_));
 sky130_fd_sc_hd__a2111o_1 _18850_ (.A1(_00303_),
    .A2(_14667_),
    .B1(_14677_),
    .C1(_14688_),
    .D1(_14706_),
    .X(_00039_));
 sky130_fd_sc_hd__nor3_1 _18851_ (.A(_12900_),
    .B(_14684_),
    .C(_12901_),
    .Y(_00040_));
 sky130_fd_sc_hd__o311ai_1 _18852_ (.A1(_12829_),
    .A2(_12836_),
    .A3(_12841_),
    .B1(is_lb_lh_lw_lbu_lhu),
    .C1(_12917_),
    .Y(_14707_));
 sky130_fd_sc_hd__nand2_1 _18853_ (.A(_13573_),
    .B(_12652_),
    .Y(_14708_));
 sky130_fd_sc_hd__a21oi_1 _18854_ (.A1(_14707_),
    .A2(_14708_),
    .B1(_14684_),
    .Y(_00044_));
 sky130_fd_sc_hd__nor2_8 _18855_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(is_slli_srli_srai),
    .Y(_01304_));
 sky130_fd_sc_hd__nand3b_2 _18856_ (.A_N(is_lui_auipc_jal),
    .B(_12855_),
    .C(_01304_),
    .Y(_14709_));
 sky130_fd_sc_hd__nor2_1 _18857_ (.A(_14709_),
    .B(_12881_),
    .Y(_14710_));
 sky130_fd_sc_hd__and4_1 _18858_ (.A(_00310_),
    .B(_12843_),
    .C(_12819_),
    .D(_00311_),
    .X(_14711_));
 sky130_fd_sc_hd__o21a_1 _18859_ (.A1(_14710_),
    .A2(_14711_),
    .B1(_14683_),
    .X(_00041_));
 sky130_fd_sc_hd__o2111ai_4 _18860_ (.A1(irq_active),
    .A2(_13540_),
    .B1(_12819_),
    .C1(_13547_),
    .D1(_13546_),
    .Y(_14712_));
 sky130_fd_sc_hd__a41oi_1 _18861_ (.A1(_12893_),
    .A2(_14712_),
    .A3(_14679_),
    .A4(_14682_),
    .B1(_12815_),
    .Y(_00038_));
 sky130_fd_sc_hd__buf_4 _18862_ (.A(_12885_),
    .X(_14713_));
 sky130_fd_sc_hd__o2111a_1 _18863_ (.A1(_14660_),
    .A2(_14669_),
    .B1(_12649_),
    .C1(_14112_),
    .D1(_14713_),
    .X(_14714_));
 sky130_fd_sc_hd__a31o_1 _18864_ (.A1(_14212_),
    .A2(_13573_),
    .A3(_14683_),
    .B1(_14714_),
    .X(_00043_));
 sky130_fd_sc_hd__buf_2 _18865_ (.A(_14696_),
    .X(_14715_));
 sky130_fd_sc_hd__buf_6 _18866_ (.A(_12670_),
    .X(_00301_));
 sky130_fd_sc_hd__a21oi_4 _18867_ (.A1(_14715_),
    .A2(_00301_),
    .B1(_13857_),
    .Y(net199));
 sky130_fd_sc_hd__nor2_8 _18868_ (.A(_00291_),
    .B(_13857_),
    .Y(net232));
 sky130_fd_sc_hd__a21o_1 _18869_ (.A1(_12635_),
    .A2(_00301_),
    .B1(_13857_),
    .X(_00316_));
 sky130_fd_sc_hd__and2_1 _18870_ (.A(_12976_),
    .B(\cpu_state[5] ),
    .X(_14716_));
 sky130_fd_sc_hd__clkbuf_1 _18871_ (.A(_14716_),
    .X(_00317_));
 sky130_fd_sc_hd__clkbuf_2 _18872_ (.A(_12845_),
    .X(_14717_));
 sky130_fd_sc_hd__buf_2 _18873_ (.A(_14717_),
    .X(_14718_));
 sky130_fd_sc_hd__nand3b_1 _18874_ (.A_N(_00307_),
    .B(_14673_),
    .C(_14689_),
    .Y(_14719_));
 sky130_fd_sc_hd__nand2_1 _18875_ (.A(_12890_),
    .B(_12816_),
    .Y(_14720_));
 sky130_fd_sc_hd__a21oi_1 _18876_ (.A1(_14702_),
    .A2(_14719_),
    .B1(_14720_),
    .Y(_14721_));
 sky130_fd_sc_hd__a21o_1 _18877_ (.A1(_12846_),
    .A2(_14683_),
    .B1(_14721_),
    .X(_14722_));
 sky130_vsdinv _18878_ (.A(_00310_),
    .Y(_14723_));
 sky130_fd_sc_hd__nor3_1 _18879_ (.A(_12811_),
    .B(_14694_),
    .C(_14720_),
    .Y(_14724_));
 sky130_fd_sc_hd__a41o_1 _18880_ (.A1(_14723_),
    .A2(_12884_),
    .A3(_12843_),
    .A4(_14699_),
    .B1(_14724_),
    .X(_14725_));
 sky130_fd_sc_hd__o32ai_4 _18881_ (.A1(_14678_),
    .A2(_14669_),
    .A3(_14640_),
    .B1(_14641_),
    .B2(_14684_),
    .Y(_14726_));
 sky130_fd_sc_hd__a221o_1 _18882_ (.A1(_14718_),
    .A2(_14722_),
    .B1(_14657_),
    .B2(_14725_),
    .C1(_14726_),
    .X(_00042_));
 sky130_fd_sc_hd__xor2_2 _18883_ (.A(_13839_),
    .B(_14266_),
    .X(_02591_));
 sky130_fd_sc_hd__nor2_4 _18884_ (.A(net354),
    .B(_14229_),
    .Y(_14727_));
 sky130_fd_sc_hd__and2_1 _18885_ (.A(net354),
    .B(_14228_),
    .X(_14728_));
 sky130_fd_sc_hd__nor2_1 _18886_ (.A(net355),
    .B(_14225_),
    .Y(_14729_));
 sky130_fd_sc_hd__and2_1 _18887_ (.A(net355),
    .B(net323),
    .X(_14730_));
 sky130_fd_sc_hd__nor2_2 _18888_ (.A(_14729_),
    .B(_14730_),
    .Y(_14731_));
 sky130_fd_sc_hd__nor2_1 _18889_ (.A(net356),
    .B(net324),
    .Y(_14732_));
 sky130_fd_sc_hd__and2_1 _18890_ (.A(net356),
    .B(net324),
    .X(_14733_));
 sky130_fd_sc_hd__nor2_2 _18891_ (.A(_14732_),
    .B(_14733_),
    .Y(_14734_));
 sky130_fd_sc_hd__nor2_1 _18892_ (.A(_13800_),
    .B(_14221_),
    .Y(_14735_));
 sky130_fd_sc_hd__and2_1 _18893_ (.A(net357),
    .B(net325),
    .X(_14736_));
 sky130_fd_sc_hd__nor2_2 _18894_ (.A(_14735_),
    .B(_14736_),
    .Y(_14737_));
 sky130_fd_sc_hd__nor3_2 _18895_ (.A(_14731_),
    .B(_14734_),
    .C(_14737_),
    .Y(_14738_));
 sky130_fd_sc_hd__nor2_1 _18896_ (.A(net359),
    .B(net327),
    .Y(_14739_));
 sky130_fd_sc_hd__and2_1 _18897_ (.A(net359),
    .B(net327),
    .X(_14740_));
 sky130_fd_sc_hd__nor2_1 _18898_ (.A(net358),
    .B(net326),
    .Y(_14741_));
 sky130_fd_sc_hd__and2_1 _18899_ (.A(net358),
    .B(net326),
    .X(_14742_));
 sky130_fd_sc_hd__nor2_4 _18900_ (.A(_13797_),
    .B(net329),
    .Y(_14743_));
 sky130_fd_sc_hd__and2_1 _18901_ (.A(net361),
    .B(net329),
    .X(_14744_));
 sky130_fd_sc_hd__or2_1 _18902_ (.A(net330),
    .B(net362),
    .X(_14745_));
 sky130_fd_sc_hd__nand2_1 _18903_ (.A(net330),
    .B(net362),
    .Y(_14746_));
 sky130_fd_sc_hd__a2bb2oi_2 _18904_ (.A1_N(_14743_),
    .A2_N(_14744_),
    .B1(_14745_),
    .B2(_14746_),
    .Y(_14747_));
 sky130_fd_sc_hd__o221a_1 _18905_ (.A1(_14739_),
    .A2(_14740_),
    .B1(_14741_),
    .B2(_14742_),
    .C1(_14747_),
    .X(_14748_));
 sky130_fd_sc_hd__o211a_1 _18906_ (.A1(_14727_),
    .A2(_14728_),
    .B1(_14738_),
    .C1(_14748_),
    .X(_14749_));
 sky130_fd_sc_hd__and2_1 _18907_ (.A(net347),
    .B(_14236_),
    .X(_14750_));
 sky130_vsdinv _18908_ (.A(_14750_),
    .Y(_14751_));
 sky130_fd_sc_hd__nor2_1 _18909_ (.A(_13812_),
    .B(_14236_),
    .Y(_14752_));
 sky130_vsdinv _18910_ (.A(_14752_),
    .Y(_14753_));
 sky130_fd_sc_hd__nor2_1 _18911_ (.A(net346),
    .B(_14238_),
    .Y(_14754_));
 sky130_fd_sc_hd__and2_1 _18912_ (.A(net346),
    .B(_14237_),
    .X(_14755_));
 sky130_fd_sc_hd__nor2_2 _18913_ (.A(_14754_),
    .B(_14755_),
    .Y(_14756_));
 sky130_fd_sc_hd__xor2_2 _18914_ (.A(net345),
    .B(_14239_),
    .X(_14757_));
 sky130_fd_sc_hd__xor2_4 _18915_ (.A(net352),
    .B(_14231_),
    .X(_14758_));
 sky130_fd_sc_hd__a2111oi_2 _18916_ (.A1(_14751_),
    .A2(_14753_),
    .B1(_14756_),
    .C1(_14757_),
    .D1(_14758_),
    .Y(_14759_));
 sky130_fd_sc_hd__nor2_2 _18917_ (.A(net350),
    .B(_14233_),
    .Y(_14760_));
 sky130_fd_sc_hd__and2_1 _18918_ (.A(net350),
    .B(_14233_),
    .X(_14761_));
 sky130_fd_sc_hd__nor2_4 _18919_ (.A(_14760_),
    .B(_14761_),
    .Y(_14762_));
 sky130_fd_sc_hd__nor2_2 _18920_ (.A(net351),
    .B(_14232_),
    .Y(_14763_));
 sky130_fd_sc_hd__and2_1 _18921_ (.A(net351),
    .B(net319),
    .X(_14764_));
 sky130_fd_sc_hd__nor2_4 _18922_ (.A(_14763_),
    .B(_14764_),
    .Y(_14765_));
 sky130_fd_sc_hd__nor2_2 _18923_ (.A(net348),
    .B(_14234_),
    .Y(_14766_));
 sky130_fd_sc_hd__and2_1 _18924_ (.A(net348),
    .B(net316),
    .X(_14767_));
 sky130_fd_sc_hd__nor2_4 _18925_ (.A(net353),
    .B(_14230_),
    .Y(_14768_));
 sky130_fd_sc_hd__and2_1 _18926_ (.A(net353),
    .B(net321),
    .X(_14769_));
 sky130_fd_sc_hd__o22ai_4 _18927_ (.A1(_14766_),
    .A2(_14767_),
    .B1(_14768_),
    .B2(_14769_),
    .Y(_14770_));
 sky130_fd_sc_hd__nor3_4 _18928_ (.A(_14762_),
    .B(_14765_),
    .C(_14770_),
    .Y(_14771_));
 sky130_fd_sc_hd__and3_1 _18929_ (.A(_14749_),
    .B(_14759_),
    .C(_14771_),
    .X(_14772_));
 sky130_vsdinv _18930_ (.A(_14772_),
    .Y(_14773_));
 sky130_fd_sc_hd__nor2_4 _18931_ (.A(_13837_),
    .B(_14263_),
    .Y(_14774_));
 sky130_fd_sc_hd__and2_1 _18932_ (.A(net492),
    .B(_14263_),
    .X(_14775_));
 sky130_fd_sc_hd__nor2_1 _18933_ (.A(_13829_),
    .B(_14257_),
    .Y(_14776_));
 sky130_fd_sc_hd__and2_1 _18934_ (.A(net227),
    .B(net333),
    .X(_14777_));
 sky130_fd_sc_hd__o22a_1 _18935_ (.A1(_14774_),
    .A2(_14775_),
    .B1(_14776_),
    .B2(_14777_),
    .X(_14778_));
 sky130_fd_sc_hd__nor2_1 _18936_ (.A(_13833_),
    .B(_14260_),
    .Y(_14779_));
 sky130_fd_sc_hd__and2_1 _18937_ (.A(_13833_),
    .B(net331),
    .X(_14780_));
 sky130_fd_sc_hd__nor2_1 _18938_ (.A(_14779_),
    .B(_14780_),
    .Y(_14781_));
 sky130_vsdinv _18939_ (.A(_14781_),
    .Y(_14782_));
 sky130_fd_sc_hd__nand3b_1 _18940_ (.A_N(_02591_),
    .B(_14778_),
    .C(_14782_),
    .Y(_14783_));
 sky130_fd_sc_hd__nor2_1 _18941_ (.A(_13825_),
    .B(_14253_),
    .Y(_14784_));
 sky130_fd_sc_hd__and2_1 _18942_ (.A(_13825_),
    .B(_14252_),
    .X(_14785_));
 sky130_fd_sc_hd__nor2_2 _18943_ (.A(_14784_),
    .B(_14785_),
    .Y(_14786_));
 sky130_fd_sc_hd__xor2_2 _18944_ (.A(_13835_),
    .B(_14261_),
    .X(_14787_));
 sky130_fd_sc_hd__nor2_1 _18945_ (.A(_13827_),
    .B(_14255_),
    .Y(_14788_));
 sky130_fd_sc_hd__and2_1 _18946_ (.A(_13827_),
    .B(_14255_),
    .X(_14789_));
 sky130_fd_sc_hd__nor2_2 _18947_ (.A(_14788_),
    .B(_14789_),
    .Y(_14790_));
 sky130_fd_sc_hd__xor2_2 _18948_ (.A(net226),
    .B(_14258_),
    .X(_14791_));
 sky130_fd_sc_hd__or4_4 _18949_ (.A(_14786_),
    .B(_14787_),
    .C(_14790_),
    .D(_14791_),
    .X(_14792_));
 sky130_fd_sc_hd__xor2_2 _18950_ (.A(net339),
    .B(_14247_),
    .X(_14793_));
 sky130_fd_sc_hd__nor2_2 _18951_ (.A(net369),
    .B(_14249_),
    .Y(_14794_));
 sky130_fd_sc_hd__and2_1 _18952_ (.A(net369),
    .B(_14249_),
    .X(_14795_));
 sky130_fd_sc_hd__nor2_1 _18953_ (.A(_14794_),
    .B(_14795_),
    .Y(_14796_));
 sky130_fd_sc_hd__xor2_2 _18954_ (.A(net368),
    .B(_14250_),
    .X(_14797_));
 sky130_fd_sc_hd__xor2_4 _18955_ (.A(net340),
    .B(_14246_),
    .X(_14798_));
 sky130_fd_sc_hd__or4_4 _18956_ (.A(_14793_),
    .B(_14796_),
    .C(_14797_),
    .D(_14798_),
    .X(_14799_));
 sky130_fd_sc_hd__nor2_2 _18957_ (.A(net343),
    .B(_14242_),
    .Y(_14800_));
 sky130_fd_sc_hd__and2_1 _18958_ (.A(net343),
    .B(net311),
    .X(_14801_));
 sky130_fd_sc_hd__nor2_4 _18959_ (.A(_14800_),
    .B(_14801_),
    .Y(_14802_));
 sky130_fd_sc_hd__nor2_2 _18960_ (.A(net344),
    .B(_14241_),
    .Y(_14803_));
 sky130_fd_sc_hd__and2_1 _18961_ (.A(net344),
    .B(net312),
    .X(_14804_));
 sky130_fd_sc_hd__nor2_4 _18962_ (.A(_14803_),
    .B(_14804_),
    .Y(_14805_));
 sky130_fd_sc_hd__nor2_4 _18963_ (.A(net342),
    .B(_14243_),
    .Y(_14806_));
 sky130_fd_sc_hd__and2_1 _18964_ (.A(net342),
    .B(net310),
    .X(_14807_));
 sky130_fd_sc_hd__nor2_8 _18965_ (.A(net341),
    .B(_14245_),
    .Y(_14808_));
 sky130_fd_sc_hd__and2_2 _18966_ (.A(net341),
    .B(_14245_),
    .X(_14809_));
 sky130_fd_sc_hd__o22ai_4 _18967_ (.A1(_14806_),
    .A2(_14807_),
    .B1(_14808_),
    .B2(_14809_),
    .Y(_14810_));
 sky130_fd_sc_hd__nor3_4 _18968_ (.A(_14802_),
    .B(_14805_),
    .C(_14810_),
    .Y(_14811_));
 sky130_fd_sc_hd__or4b_4 _18969_ (.A(_14783_),
    .B(_14792_),
    .C(_14799_),
    .D_N(_14811_),
    .X(_14812_));
 sky130_fd_sc_hd__nor2_4 _18970_ (.A(_14773_),
    .B(_14812_),
    .Y(_00000_));
 sky130_fd_sc_hd__a21oi_1 _18971_ (.A1(_12799_),
    .A2(_12801_),
    .B1(_12791_),
    .Y(\pcpi_mul.instr_any_mulh ));
 sky130_fd_sc_hd__nand2b_1 _18972_ (.A_N(instr_blt),
    .B(_13570_),
    .Y(_00006_));
 sky130_fd_sc_hd__nand2b_1 _18973_ (.A_N(instr_bltu),
    .B(_13569_),
    .Y(_00007_));
 sky130_fd_sc_hd__o21ai_1 _18974_ (.A1(_12633_),
    .A2(_12634_),
    .B1(_12676_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand3b_1 _18975_ (.A_N(_12976_),
    .B(_12648_),
    .C(_14212_),
    .Y(_14813_));
 sky130_vsdinv _18976_ (.A(_14813_),
    .Y(_14814_));
 sky130_fd_sc_hd__a21oi_1 _18977_ (.A1(_14195_),
    .A2(_12657_),
    .B1(_13093_),
    .Y(_14815_));
 sky130_fd_sc_hd__a21oi_1 _18978_ (.A1(instr_sh),
    .A2(_14814_),
    .B1(_14815_),
    .Y(_14816_));
 sky130_vsdinv _18979_ (.A(_14658_),
    .Y(_14817_));
 sky130_fd_sc_hd__clkbuf_2 _18980_ (.A(_14817_),
    .X(_14818_));
 sky130_fd_sc_hd__a2bb2oi_1 _18981_ (.A1_N(_00319_),
    .A2_N(_00317_),
    .B1(_12640_),
    .B2(_12639_),
    .Y(_14819_));
 sky130_fd_sc_hd__o211a_1 _18982_ (.A1(_12651_),
    .A2(_14212_),
    .B1(_12640_),
    .C1(_12890_),
    .X(_14820_));
 sky130_fd_sc_hd__a2111oi_2 _18983_ (.A1(_12848_),
    .A2(_00297_),
    .B1(_12642_),
    .C1(_14819_),
    .D1(_14820_),
    .Y(_14821_));
 sky130_fd_sc_hd__o22ai_1 _18984_ (.A1(_00296_),
    .A2(_14816_),
    .B1(_14818_),
    .B2(_14821_),
    .Y(_00047_));
 sky130_fd_sc_hd__clkbuf_4 _18985_ (.A(_14717_),
    .X(_14822_));
 sky130_fd_sc_hd__nor3_2 _18986_ (.A(_14822_),
    .B(_12652_),
    .C(_14212_),
    .Y(_00336_));
 sky130_fd_sc_hd__o2111ai_4 _18987_ (.A1(_12666_),
    .A2(_13089_),
    .B1(_12650_),
    .C1(net456),
    .D1(_12632_),
    .Y(_00338_));
 sky130_vsdinv _18988_ (.A(alu_eq),
    .Y(_00340_));
 sky130_fd_sc_hd__nor3_2 _18989_ (.A(instr_bne),
    .B(is_slti_blt_slt),
    .C(is_sltiu_bltu_sltu),
    .Y(_14823_));
 sky130_fd_sc_hd__nor3b_4 _18990_ (.A(instr_bgeu),
    .B(instr_bge),
    .C_N(_14823_),
    .Y(_00341_));
 sky130_fd_sc_hd__and2b_1 _18991_ (.A_N(alu_ltu),
    .B(instr_bgeu),
    .X(_14824_));
 sky130_fd_sc_hd__and2b_1 _18992_ (.A_N(alu_lts),
    .B(instr_bge),
    .X(_14825_));
 sky130_fd_sc_hd__a221o_1 _18993_ (.A1(_00340_),
    .A2(instr_bne),
    .B1(is_slti_blt_slt),
    .B2(alu_lts),
    .C1(_14825_),
    .X(_14826_));
 sky130_fd_sc_hd__a211oi_4 _18994_ (.A1(is_sltiu_bltu_sltu),
    .A2(alu_ltu),
    .B1(_14824_),
    .C1(_14826_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand3b_1 _18995_ (.A_N(_12639_),
    .B(_12666_),
    .C(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__o22ai_1 _18996_ (.A1(_00346_),
    .A2(_12813_),
    .B1(_00339_),
    .B2(_00297_),
    .Y(_00347_));
 sky130_fd_sc_hd__o21ba_1 _18997_ (.A1(_13048_),
    .A2(do_waitirq),
    .B1_N(_12863_),
    .X(_00349_));
 sky130_fd_sc_hd__nor3b_1 _18998_ (.A(_13558_),
    .B(_13564_),
    .C_N(_00349_),
    .Y(_00351_));
 sky130_fd_sc_hd__buf_2 _18999_ (.A(_12885_),
    .X(_14827_));
 sky130_fd_sc_hd__nor3_2 _19000_ (.A(_14822_),
    .B(_12917_),
    .C(_14827_),
    .Y(_00354_));
 sky130_fd_sc_hd__a211oi_1 _19001_ (.A1(_14822_),
    .A2(_12640_),
    .B1(_12917_),
    .C1(_14827_),
    .Y(_00355_));
 sky130_vsdinv _19002_ (.A(\cpuregs[0][1] ),
    .Y(_00371_));
 sky130_vsdinv _19003_ (.A(\cpuregs[1][1] ),
    .Y(_00372_));
 sky130_vsdinv _19004_ (.A(\cpuregs[2][1] ),
    .Y(_00373_));
 sky130_vsdinv _19005_ (.A(\cpuregs[3][1] ),
    .Y(_00374_));
 sky130_vsdinv _19006_ (.A(\cpuregs[4][1] ),
    .Y(_00376_));
 sky130_vsdinv _19007_ (.A(\cpuregs[5][1] ),
    .Y(_00377_));
 sky130_vsdinv _19008_ (.A(\cpuregs[6][1] ),
    .Y(_00378_));
 sky130_vsdinv _19009_ (.A(\cpuregs[7][1] ),
    .Y(_00379_));
 sky130_vsdinv _19010_ (.A(\cpuregs[8][1] ),
    .Y(_00381_));
 sky130_vsdinv _19011_ (.A(\cpuregs[9][1] ),
    .Y(_00382_));
 sky130_vsdinv _19012_ (.A(\cpuregs[10][1] ),
    .Y(_00383_));
 sky130_vsdinv _19013_ (.A(\cpuregs[11][1] ),
    .Y(_00384_));
 sky130_vsdinv _19014_ (.A(\cpuregs[12][1] ),
    .Y(_00386_));
 sky130_vsdinv _19015_ (.A(\cpuregs[13][1] ),
    .Y(_00387_));
 sky130_vsdinv _19016_ (.A(\cpuregs[14][1] ),
    .Y(_00388_));
 sky130_vsdinv _19017_ (.A(\cpuregs[15][1] ),
    .Y(_00389_));
 sky130_vsdinv _19018_ (.A(\cpuregs[16][1] ),
    .Y(_00392_));
 sky130_vsdinv _19019_ (.A(\cpuregs[17][1] ),
    .Y(_00393_));
 sky130_vsdinv _19020_ (.A(\cpuregs[18][1] ),
    .Y(_00394_));
 sky130_vsdinv _19021_ (.A(\cpuregs[19][1] ),
    .Y(_00395_));
 sky130_vsdinv _19022_ (.A(_12846_),
    .Y(_00302_));
 sky130_vsdinv _19023_ (.A(\cpuregs[0][2] ),
    .Y(_00398_));
 sky130_vsdinv _19024_ (.A(\cpuregs[1][2] ),
    .Y(_00399_));
 sky130_vsdinv _19025_ (.A(\cpuregs[2][2] ),
    .Y(_00400_));
 sky130_vsdinv _19026_ (.A(\cpuregs[3][2] ),
    .Y(_00401_));
 sky130_vsdinv _19027_ (.A(\cpuregs[4][2] ),
    .Y(_00403_));
 sky130_vsdinv _19028_ (.A(\cpuregs[5][2] ),
    .Y(_00404_));
 sky130_vsdinv _19029_ (.A(\cpuregs[6][2] ),
    .Y(_00405_));
 sky130_vsdinv _19030_ (.A(\cpuregs[7][2] ),
    .Y(_00406_));
 sky130_vsdinv _19031_ (.A(\cpuregs[8][2] ),
    .Y(_00408_));
 sky130_vsdinv _19032_ (.A(\cpuregs[9][2] ),
    .Y(_00409_));
 sky130_vsdinv _19033_ (.A(\cpuregs[10][2] ),
    .Y(_00410_));
 sky130_vsdinv _19034_ (.A(\cpuregs[11][2] ),
    .Y(_00411_));
 sky130_vsdinv _19035_ (.A(\cpuregs[12][2] ),
    .Y(_00413_));
 sky130_vsdinv _19036_ (.A(\cpuregs[13][2] ),
    .Y(_00414_));
 sky130_vsdinv _19037_ (.A(\cpuregs[14][2] ),
    .Y(_00415_));
 sky130_vsdinv _19038_ (.A(\cpuregs[15][2] ),
    .Y(_00416_));
 sky130_vsdinv _19039_ (.A(\cpuregs[16][2] ),
    .Y(_00419_));
 sky130_vsdinv _19040_ (.A(\cpuregs[17][2] ),
    .Y(_00420_));
 sky130_vsdinv _19041_ (.A(\cpuregs[18][2] ),
    .Y(_00421_));
 sky130_vsdinv _19042_ (.A(\cpuregs[19][2] ),
    .Y(_00422_));
 sky130_vsdinv _19043_ (.A(\cpuregs[0][3] ),
    .Y(_00425_));
 sky130_vsdinv _19044_ (.A(\cpuregs[1][3] ),
    .Y(_00426_));
 sky130_vsdinv _19045_ (.A(\cpuregs[2][3] ),
    .Y(_00427_));
 sky130_vsdinv _19046_ (.A(\cpuregs[3][3] ),
    .Y(_00428_));
 sky130_vsdinv _19047_ (.A(\cpuregs[4][3] ),
    .Y(_00430_));
 sky130_vsdinv _19048_ (.A(\cpuregs[5][3] ),
    .Y(_00431_));
 sky130_vsdinv _19049_ (.A(\cpuregs[6][3] ),
    .Y(_00432_));
 sky130_vsdinv _19050_ (.A(\cpuregs[7][3] ),
    .Y(_00433_));
 sky130_vsdinv _19051_ (.A(\cpuregs[8][3] ),
    .Y(_00435_));
 sky130_vsdinv _19052_ (.A(\cpuregs[9][3] ),
    .Y(_00436_));
 sky130_vsdinv _19053_ (.A(\cpuregs[10][3] ),
    .Y(_00437_));
 sky130_vsdinv _19054_ (.A(\cpuregs[11][3] ),
    .Y(_00438_));
 sky130_vsdinv _19055_ (.A(\cpuregs[12][3] ),
    .Y(_00440_));
 sky130_vsdinv _19056_ (.A(\cpuregs[13][3] ),
    .Y(_00441_));
 sky130_vsdinv _19057_ (.A(\cpuregs[14][3] ),
    .Y(_00442_));
 sky130_vsdinv _19058_ (.A(\cpuregs[15][3] ),
    .Y(_00443_));
 sky130_vsdinv _19059_ (.A(\cpuregs[16][3] ),
    .Y(_00446_));
 sky130_vsdinv _19060_ (.A(\cpuregs[17][3] ),
    .Y(_00447_));
 sky130_vsdinv _19061_ (.A(\cpuregs[18][3] ),
    .Y(_00448_));
 sky130_vsdinv _19062_ (.A(\cpuregs[19][3] ),
    .Y(_00449_));
 sky130_vsdinv _19063_ (.A(\cpuregs[0][4] ),
    .Y(_00452_));
 sky130_vsdinv _19064_ (.A(\cpuregs[1][4] ),
    .Y(_00453_));
 sky130_vsdinv _19065_ (.A(\cpuregs[2][4] ),
    .Y(_00454_));
 sky130_vsdinv _19066_ (.A(\cpuregs[3][4] ),
    .Y(_00455_));
 sky130_vsdinv _19067_ (.A(\cpuregs[4][4] ),
    .Y(_00457_));
 sky130_vsdinv _19068_ (.A(\cpuregs[5][4] ),
    .Y(_00458_));
 sky130_vsdinv _19069_ (.A(\cpuregs[6][4] ),
    .Y(_00459_));
 sky130_vsdinv _19070_ (.A(\cpuregs[7][4] ),
    .Y(_00460_));
 sky130_vsdinv _19071_ (.A(\cpuregs[8][4] ),
    .Y(_00462_));
 sky130_vsdinv _19072_ (.A(\cpuregs[9][4] ),
    .Y(_00463_));
 sky130_vsdinv _19073_ (.A(\cpuregs[10][4] ),
    .Y(_00464_));
 sky130_vsdinv _19074_ (.A(\cpuregs[11][4] ),
    .Y(_00465_));
 sky130_vsdinv _19075_ (.A(\cpuregs[12][4] ),
    .Y(_00467_));
 sky130_vsdinv _19076_ (.A(\cpuregs[13][4] ),
    .Y(_00468_));
 sky130_vsdinv _19077_ (.A(\cpuregs[14][4] ),
    .Y(_00469_));
 sky130_vsdinv _19078_ (.A(\cpuregs[15][4] ),
    .Y(_00470_));
 sky130_vsdinv _19079_ (.A(\cpuregs[16][4] ),
    .Y(_00473_));
 sky130_vsdinv _19080_ (.A(\cpuregs[17][4] ),
    .Y(_00474_));
 sky130_vsdinv _19081_ (.A(\cpuregs[18][4] ),
    .Y(_00475_));
 sky130_vsdinv _19082_ (.A(\cpuregs[19][4] ),
    .Y(_00476_));
 sky130_vsdinv _19083_ (.A(\cpuregs[0][5] ),
    .Y(_00479_));
 sky130_vsdinv _19084_ (.A(\cpuregs[1][5] ),
    .Y(_00480_));
 sky130_vsdinv _19085_ (.A(\cpuregs[2][5] ),
    .Y(_00481_));
 sky130_vsdinv _19086_ (.A(\cpuregs[3][5] ),
    .Y(_00482_));
 sky130_vsdinv _19087_ (.A(\cpuregs[4][5] ),
    .Y(_00484_));
 sky130_vsdinv _19088_ (.A(\cpuregs[5][5] ),
    .Y(_00485_));
 sky130_vsdinv _19089_ (.A(\cpuregs[6][5] ),
    .Y(_00486_));
 sky130_vsdinv _19090_ (.A(\cpuregs[7][5] ),
    .Y(_00487_));
 sky130_vsdinv _19091_ (.A(\cpuregs[8][5] ),
    .Y(_00489_));
 sky130_vsdinv _19092_ (.A(\cpuregs[9][5] ),
    .Y(_00490_));
 sky130_vsdinv _19093_ (.A(\cpuregs[10][5] ),
    .Y(_00491_));
 sky130_vsdinv _19094_ (.A(\cpuregs[11][5] ),
    .Y(_00492_));
 sky130_vsdinv _19095_ (.A(\cpuregs[12][5] ),
    .Y(_00494_));
 sky130_vsdinv _19096_ (.A(\cpuregs[13][5] ),
    .Y(_00495_));
 sky130_vsdinv _19097_ (.A(\cpuregs[14][5] ),
    .Y(_00496_));
 sky130_vsdinv _19098_ (.A(\cpuregs[15][5] ),
    .Y(_00497_));
 sky130_vsdinv _19099_ (.A(\cpuregs[16][5] ),
    .Y(_00500_));
 sky130_vsdinv _19100_ (.A(\cpuregs[17][5] ),
    .Y(_00501_));
 sky130_vsdinv _19101_ (.A(\cpuregs[18][5] ),
    .Y(_00502_));
 sky130_vsdinv _19102_ (.A(\cpuregs[19][5] ),
    .Y(_00503_));
 sky130_vsdinv _19103_ (.A(\cpuregs[0][6] ),
    .Y(_00506_));
 sky130_vsdinv _19104_ (.A(\cpuregs[1][6] ),
    .Y(_00507_));
 sky130_vsdinv _19105_ (.A(\cpuregs[2][6] ),
    .Y(_00508_));
 sky130_vsdinv _19106_ (.A(\cpuregs[3][6] ),
    .Y(_00509_));
 sky130_vsdinv _19107_ (.A(\cpuregs[4][6] ),
    .Y(_00511_));
 sky130_vsdinv _19108_ (.A(\cpuregs[5][6] ),
    .Y(_00512_));
 sky130_vsdinv _19109_ (.A(\cpuregs[6][6] ),
    .Y(_00513_));
 sky130_vsdinv _19110_ (.A(\cpuregs[7][6] ),
    .Y(_00514_));
 sky130_vsdinv _19111_ (.A(\cpuregs[8][6] ),
    .Y(_00516_));
 sky130_vsdinv _19112_ (.A(\cpuregs[9][6] ),
    .Y(_00517_));
 sky130_vsdinv _19113_ (.A(\cpuregs[10][6] ),
    .Y(_00518_));
 sky130_vsdinv _19114_ (.A(\cpuregs[11][6] ),
    .Y(_00519_));
 sky130_vsdinv _19115_ (.A(\cpuregs[12][6] ),
    .Y(_00521_));
 sky130_vsdinv _19116_ (.A(\cpuregs[13][6] ),
    .Y(_00522_));
 sky130_vsdinv _19117_ (.A(\cpuregs[14][6] ),
    .Y(_00523_));
 sky130_vsdinv _19118_ (.A(\cpuregs[15][6] ),
    .Y(_00524_));
 sky130_vsdinv _19119_ (.A(\cpuregs[16][6] ),
    .Y(_00527_));
 sky130_vsdinv _19120_ (.A(\cpuregs[17][6] ),
    .Y(_00528_));
 sky130_vsdinv _19121_ (.A(\cpuregs[18][6] ),
    .Y(_00529_));
 sky130_vsdinv _19122_ (.A(\cpuregs[19][6] ),
    .Y(_00530_));
 sky130_vsdinv _19123_ (.A(\cpuregs[0][7] ),
    .Y(_00533_));
 sky130_vsdinv _19124_ (.A(\cpuregs[1][7] ),
    .Y(_00534_));
 sky130_vsdinv _19125_ (.A(\cpuregs[2][7] ),
    .Y(_00535_));
 sky130_vsdinv _19126_ (.A(\cpuregs[3][7] ),
    .Y(_00536_));
 sky130_vsdinv _19127_ (.A(\cpuregs[4][7] ),
    .Y(_00538_));
 sky130_vsdinv _19128_ (.A(\cpuregs[5][7] ),
    .Y(_00539_));
 sky130_vsdinv _19129_ (.A(\cpuregs[6][7] ),
    .Y(_00540_));
 sky130_vsdinv _19130_ (.A(\cpuregs[7][7] ),
    .Y(_00541_));
 sky130_vsdinv _19131_ (.A(\cpuregs[8][7] ),
    .Y(_00543_));
 sky130_vsdinv _19132_ (.A(\cpuregs[9][7] ),
    .Y(_00544_));
 sky130_vsdinv _19133_ (.A(\cpuregs[10][7] ),
    .Y(_00545_));
 sky130_vsdinv _19134_ (.A(\cpuregs[11][7] ),
    .Y(_00546_));
 sky130_vsdinv _19135_ (.A(\cpuregs[12][7] ),
    .Y(_00548_));
 sky130_vsdinv _19136_ (.A(\cpuregs[13][7] ),
    .Y(_00549_));
 sky130_vsdinv _19137_ (.A(\cpuregs[14][7] ),
    .Y(_00550_));
 sky130_vsdinv _19138_ (.A(\cpuregs[15][7] ),
    .Y(_00551_));
 sky130_vsdinv _19139_ (.A(\cpuregs[16][7] ),
    .Y(_00554_));
 sky130_vsdinv _19140_ (.A(\cpuregs[17][7] ),
    .Y(_00555_));
 sky130_vsdinv _19141_ (.A(\cpuregs[18][7] ),
    .Y(_00556_));
 sky130_vsdinv _19142_ (.A(\cpuregs[19][7] ),
    .Y(_00557_));
 sky130_vsdinv _19143_ (.A(\cpuregs[0][8] ),
    .Y(_00560_));
 sky130_vsdinv _19144_ (.A(\cpuregs[1][8] ),
    .Y(_00561_));
 sky130_vsdinv _19145_ (.A(\cpuregs[2][8] ),
    .Y(_00562_));
 sky130_vsdinv _19146_ (.A(\cpuregs[3][8] ),
    .Y(_00563_));
 sky130_vsdinv _19147_ (.A(\cpuregs[4][8] ),
    .Y(_00565_));
 sky130_vsdinv _19148_ (.A(\cpuregs[5][8] ),
    .Y(_00566_));
 sky130_vsdinv _19149_ (.A(\cpuregs[6][8] ),
    .Y(_00567_));
 sky130_vsdinv _19150_ (.A(\cpuregs[7][8] ),
    .Y(_00568_));
 sky130_vsdinv _19151_ (.A(\cpuregs[8][8] ),
    .Y(_00570_));
 sky130_vsdinv _19152_ (.A(\cpuregs[9][8] ),
    .Y(_00571_));
 sky130_vsdinv _19153_ (.A(\cpuregs[10][8] ),
    .Y(_00572_));
 sky130_vsdinv _19154_ (.A(\cpuregs[11][8] ),
    .Y(_00573_));
 sky130_vsdinv _19155_ (.A(\cpuregs[12][8] ),
    .Y(_00575_));
 sky130_vsdinv _19156_ (.A(\cpuregs[13][8] ),
    .Y(_00576_));
 sky130_vsdinv _19157_ (.A(\cpuregs[14][8] ),
    .Y(_00577_));
 sky130_vsdinv _19158_ (.A(\cpuregs[15][8] ),
    .Y(_00578_));
 sky130_vsdinv _19159_ (.A(\cpuregs[16][8] ),
    .Y(_00581_));
 sky130_vsdinv _19160_ (.A(\cpuregs[17][8] ),
    .Y(_00582_));
 sky130_vsdinv _19161_ (.A(\cpuregs[18][8] ),
    .Y(_00583_));
 sky130_vsdinv _19162_ (.A(\cpuregs[19][8] ),
    .Y(_00584_));
 sky130_vsdinv _19163_ (.A(\cpuregs[0][9] ),
    .Y(_00587_));
 sky130_vsdinv _19164_ (.A(\cpuregs[1][9] ),
    .Y(_00588_));
 sky130_vsdinv _19165_ (.A(\cpuregs[2][9] ),
    .Y(_00589_));
 sky130_vsdinv _19166_ (.A(\cpuregs[3][9] ),
    .Y(_00590_));
 sky130_vsdinv _19167_ (.A(\cpuregs[4][9] ),
    .Y(_00592_));
 sky130_vsdinv _19168_ (.A(\cpuregs[5][9] ),
    .Y(_00593_));
 sky130_vsdinv _19169_ (.A(\cpuregs[6][9] ),
    .Y(_00594_));
 sky130_vsdinv _19170_ (.A(\cpuregs[7][9] ),
    .Y(_00595_));
 sky130_vsdinv _19171_ (.A(\cpuregs[8][9] ),
    .Y(_00597_));
 sky130_vsdinv _19172_ (.A(\cpuregs[9][9] ),
    .Y(_00598_));
 sky130_vsdinv _19173_ (.A(\cpuregs[10][9] ),
    .Y(_00599_));
 sky130_vsdinv _19174_ (.A(\cpuregs[11][9] ),
    .Y(_00600_));
 sky130_vsdinv _19175_ (.A(\cpuregs[12][9] ),
    .Y(_00602_));
 sky130_vsdinv _19176_ (.A(\cpuregs[13][9] ),
    .Y(_00603_));
 sky130_vsdinv _19177_ (.A(\cpuregs[14][9] ),
    .Y(_00604_));
 sky130_vsdinv _19178_ (.A(\cpuregs[15][9] ),
    .Y(_00605_));
 sky130_vsdinv _19179_ (.A(\cpuregs[16][9] ),
    .Y(_00608_));
 sky130_vsdinv _19180_ (.A(\cpuregs[17][9] ),
    .Y(_00609_));
 sky130_vsdinv _19181_ (.A(\cpuregs[18][9] ),
    .Y(_00610_));
 sky130_vsdinv _19182_ (.A(\cpuregs[19][9] ),
    .Y(_00611_));
 sky130_vsdinv _19183_ (.A(\cpuregs[0][10] ),
    .Y(_00614_));
 sky130_vsdinv _19184_ (.A(\cpuregs[1][10] ),
    .Y(_00615_));
 sky130_vsdinv _19185_ (.A(\cpuregs[2][10] ),
    .Y(_00616_));
 sky130_vsdinv _19186_ (.A(\cpuregs[3][10] ),
    .Y(_00617_));
 sky130_vsdinv _19187_ (.A(\cpuregs[4][10] ),
    .Y(_00619_));
 sky130_vsdinv _19188_ (.A(\cpuregs[5][10] ),
    .Y(_00620_));
 sky130_vsdinv _19189_ (.A(\cpuregs[6][10] ),
    .Y(_00621_));
 sky130_vsdinv _19190_ (.A(\cpuregs[7][10] ),
    .Y(_00622_));
 sky130_vsdinv _19191_ (.A(\cpuregs[8][10] ),
    .Y(_00624_));
 sky130_vsdinv _19192_ (.A(\cpuregs[9][10] ),
    .Y(_00625_));
 sky130_vsdinv _19193_ (.A(\cpuregs[10][10] ),
    .Y(_00626_));
 sky130_vsdinv _19194_ (.A(\cpuregs[11][10] ),
    .Y(_00627_));
 sky130_vsdinv _19195_ (.A(\cpuregs[12][10] ),
    .Y(_00629_));
 sky130_vsdinv _19196_ (.A(\cpuregs[13][10] ),
    .Y(_00630_));
 sky130_vsdinv _19197_ (.A(\cpuregs[14][10] ),
    .Y(_00631_));
 sky130_vsdinv _19198_ (.A(\cpuregs[15][10] ),
    .Y(_00632_));
 sky130_vsdinv _19199_ (.A(\cpuregs[16][10] ),
    .Y(_00635_));
 sky130_vsdinv _19200_ (.A(\cpuregs[17][10] ),
    .Y(_00636_));
 sky130_vsdinv _19201_ (.A(\cpuregs[18][10] ),
    .Y(_00637_));
 sky130_vsdinv _19202_ (.A(\cpuregs[19][10] ),
    .Y(_00638_));
 sky130_vsdinv _19203_ (.A(\cpuregs[0][11] ),
    .Y(_00641_));
 sky130_vsdinv _19204_ (.A(\cpuregs[1][11] ),
    .Y(_00642_));
 sky130_vsdinv _19205_ (.A(\cpuregs[2][11] ),
    .Y(_00643_));
 sky130_vsdinv _19206_ (.A(\cpuregs[3][11] ),
    .Y(_00644_));
 sky130_vsdinv _19207_ (.A(\cpuregs[4][11] ),
    .Y(_00646_));
 sky130_vsdinv _19208_ (.A(\cpuregs[5][11] ),
    .Y(_00647_));
 sky130_vsdinv _19209_ (.A(\cpuregs[6][11] ),
    .Y(_00648_));
 sky130_vsdinv _19210_ (.A(\cpuregs[7][11] ),
    .Y(_00649_));
 sky130_vsdinv _19211_ (.A(\cpuregs[8][11] ),
    .Y(_00651_));
 sky130_vsdinv _19212_ (.A(\cpuregs[9][11] ),
    .Y(_00652_));
 sky130_vsdinv _19213_ (.A(\cpuregs[10][11] ),
    .Y(_00653_));
 sky130_vsdinv _19214_ (.A(\cpuregs[11][11] ),
    .Y(_00654_));
 sky130_vsdinv _19215_ (.A(\cpuregs[12][11] ),
    .Y(_00656_));
 sky130_vsdinv _19216_ (.A(\cpuregs[13][11] ),
    .Y(_00657_));
 sky130_vsdinv _19217_ (.A(\cpuregs[14][11] ),
    .Y(_00658_));
 sky130_vsdinv _19218_ (.A(\cpuregs[15][11] ),
    .Y(_00659_));
 sky130_vsdinv _19219_ (.A(\cpuregs[16][11] ),
    .Y(_00662_));
 sky130_vsdinv _19220_ (.A(\cpuregs[17][11] ),
    .Y(_00663_));
 sky130_vsdinv _19221_ (.A(\cpuregs[18][11] ),
    .Y(_00664_));
 sky130_vsdinv _19222_ (.A(\cpuregs[19][11] ),
    .Y(_00665_));
 sky130_vsdinv _19223_ (.A(\cpuregs[0][12] ),
    .Y(_00668_));
 sky130_vsdinv _19224_ (.A(\cpuregs[1][12] ),
    .Y(_00669_));
 sky130_vsdinv _19225_ (.A(\cpuregs[2][12] ),
    .Y(_00670_));
 sky130_vsdinv _19226_ (.A(\cpuregs[3][12] ),
    .Y(_00671_));
 sky130_vsdinv _19227_ (.A(\cpuregs[4][12] ),
    .Y(_00673_));
 sky130_vsdinv _19228_ (.A(\cpuregs[5][12] ),
    .Y(_00674_));
 sky130_vsdinv _19229_ (.A(\cpuregs[6][12] ),
    .Y(_00675_));
 sky130_vsdinv _19230_ (.A(\cpuregs[7][12] ),
    .Y(_00676_));
 sky130_vsdinv _19231_ (.A(\cpuregs[8][12] ),
    .Y(_00678_));
 sky130_vsdinv _19232_ (.A(\cpuregs[9][12] ),
    .Y(_00679_));
 sky130_vsdinv _19233_ (.A(\cpuregs[10][12] ),
    .Y(_00680_));
 sky130_vsdinv _19234_ (.A(\cpuregs[11][12] ),
    .Y(_00681_));
 sky130_vsdinv _19235_ (.A(\cpuregs[12][12] ),
    .Y(_00683_));
 sky130_vsdinv _19236_ (.A(\cpuregs[13][12] ),
    .Y(_00684_));
 sky130_vsdinv _19237_ (.A(\cpuregs[14][12] ),
    .Y(_00685_));
 sky130_vsdinv _19238_ (.A(\cpuregs[15][12] ),
    .Y(_00686_));
 sky130_vsdinv _19239_ (.A(\cpuregs[16][12] ),
    .Y(_00689_));
 sky130_vsdinv _19240_ (.A(\cpuregs[17][12] ),
    .Y(_00690_));
 sky130_vsdinv _19241_ (.A(\cpuregs[18][12] ),
    .Y(_00691_));
 sky130_vsdinv _19242_ (.A(\cpuregs[19][12] ),
    .Y(_00692_));
 sky130_vsdinv _19243_ (.A(\cpuregs[0][13] ),
    .Y(_00695_));
 sky130_vsdinv _19244_ (.A(\cpuregs[1][13] ),
    .Y(_00696_));
 sky130_vsdinv _19245_ (.A(\cpuregs[2][13] ),
    .Y(_00697_));
 sky130_vsdinv _19246_ (.A(\cpuregs[3][13] ),
    .Y(_00698_));
 sky130_vsdinv _19247_ (.A(\cpuregs[4][13] ),
    .Y(_00700_));
 sky130_vsdinv _19248_ (.A(\cpuregs[5][13] ),
    .Y(_00701_));
 sky130_vsdinv _19249_ (.A(\cpuregs[6][13] ),
    .Y(_00702_));
 sky130_vsdinv _19250_ (.A(\cpuregs[7][13] ),
    .Y(_00703_));
 sky130_vsdinv _19251_ (.A(\cpuregs[8][13] ),
    .Y(_00705_));
 sky130_vsdinv _19252_ (.A(\cpuregs[9][13] ),
    .Y(_00706_));
 sky130_vsdinv _19253_ (.A(\cpuregs[10][13] ),
    .Y(_00707_));
 sky130_vsdinv _19254_ (.A(\cpuregs[11][13] ),
    .Y(_00708_));
 sky130_vsdinv _19255_ (.A(\cpuregs[12][13] ),
    .Y(_00710_));
 sky130_vsdinv _19256_ (.A(\cpuregs[13][13] ),
    .Y(_00711_));
 sky130_vsdinv _19257_ (.A(\cpuregs[14][13] ),
    .Y(_00712_));
 sky130_vsdinv _19258_ (.A(\cpuregs[15][13] ),
    .Y(_00713_));
 sky130_vsdinv _19259_ (.A(\cpuregs[16][13] ),
    .Y(_00716_));
 sky130_vsdinv _19260_ (.A(\cpuregs[17][13] ),
    .Y(_00717_));
 sky130_vsdinv _19261_ (.A(\cpuregs[18][13] ),
    .Y(_00718_));
 sky130_vsdinv _19262_ (.A(\cpuregs[19][13] ),
    .Y(_00719_));
 sky130_vsdinv _19263_ (.A(\cpuregs[0][14] ),
    .Y(_00722_));
 sky130_vsdinv _19264_ (.A(\cpuregs[1][14] ),
    .Y(_00723_));
 sky130_vsdinv _19265_ (.A(\cpuregs[2][14] ),
    .Y(_00724_));
 sky130_vsdinv _19266_ (.A(\cpuregs[3][14] ),
    .Y(_00725_));
 sky130_vsdinv _19267_ (.A(\cpuregs[4][14] ),
    .Y(_00727_));
 sky130_vsdinv _19268_ (.A(\cpuregs[5][14] ),
    .Y(_00728_));
 sky130_vsdinv _19269_ (.A(\cpuregs[6][14] ),
    .Y(_00729_));
 sky130_vsdinv _19270_ (.A(\cpuregs[7][14] ),
    .Y(_00730_));
 sky130_vsdinv _19271_ (.A(\cpuregs[8][14] ),
    .Y(_00732_));
 sky130_vsdinv _19272_ (.A(\cpuregs[9][14] ),
    .Y(_00733_));
 sky130_vsdinv _19273_ (.A(\cpuregs[10][14] ),
    .Y(_00734_));
 sky130_vsdinv _19274_ (.A(\cpuregs[11][14] ),
    .Y(_00735_));
 sky130_vsdinv _19275_ (.A(\cpuregs[12][14] ),
    .Y(_00737_));
 sky130_vsdinv _19276_ (.A(\cpuregs[13][14] ),
    .Y(_00738_));
 sky130_vsdinv _19277_ (.A(\cpuregs[14][14] ),
    .Y(_00739_));
 sky130_vsdinv _19278_ (.A(\cpuregs[15][14] ),
    .Y(_00740_));
 sky130_vsdinv _19279_ (.A(\cpuregs[16][14] ),
    .Y(_00743_));
 sky130_vsdinv _19280_ (.A(\cpuregs[17][14] ),
    .Y(_00744_));
 sky130_vsdinv _19281_ (.A(\cpuregs[18][14] ),
    .Y(_00745_));
 sky130_vsdinv _19282_ (.A(\cpuregs[19][14] ),
    .Y(_00746_));
 sky130_vsdinv _19283_ (.A(\cpuregs[0][15] ),
    .Y(_00749_));
 sky130_vsdinv _19284_ (.A(\cpuregs[1][15] ),
    .Y(_00750_));
 sky130_vsdinv _19285_ (.A(\cpuregs[2][15] ),
    .Y(_00751_));
 sky130_vsdinv _19286_ (.A(\cpuregs[3][15] ),
    .Y(_00752_));
 sky130_vsdinv _19287_ (.A(\cpuregs[4][15] ),
    .Y(_00754_));
 sky130_vsdinv _19288_ (.A(\cpuregs[5][15] ),
    .Y(_00755_));
 sky130_vsdinv _19289_ (.A(\cpuregs[6][15] ),
    .Y(_00756_));
 sky130_vsdinv _19290_ (.A(\cpuregs[7][15] ),
    .Y(_00757_));
 sky130_vsdinv _19291_ (.A(\cpuregs[8][15] ),
    .Y(_00759_));
 sky130_vsdinv _19292_ (.A(\cpuregs[9][15] ),
    .Y(_00760_));
 sky130_vsdinv _19293_ (.A(\cpuregs[10][15] ),
    .Y(_00761_));
 sky130_vsdinv _19294_ (.A(\cpuregs[11][15] ),
    .Y(_00762_));
 sky130_vsdinv _19295_ (.A(\cpuregs[12][15] ),
    .Y(_00764_));
 sky130_vsdinv _19296_ (.A(\cpuregs[13][15] ),
    .Y(_00765_));
 sky130_vsdinv _19297_ (.A(\cpuregs[14][15] ),
    .Y(_00766_));
 sky130_vsdinv _19298_ (.A(\cpuregs[15][15] ),
    .Y(_00767_));
 sky130_vsdinv _19299_ (.A(\cpuregs[16][15] ),
    .Y(_00770_));
 sky130_vsdinv _19300_ (.A(\cpuregs[17][15] ),
    .Y(_00771_));
 sky130_vsdinv _19301_ (.A(\cpuregs[18][15] ),
    .Y(_00772_));
 sky130_vsdinv _19302_ (.A(\cpuregs[19][15] ),
    .Y(_00773_));
 sky130_vsdinv _19303_ (.A(\cpuregs[0][16] ),
    .Y(_00776_));
 sky130_vsdinv _19304_ (.A(\cpuregs[1][16] ),
    .Y(_00777_));
 sky130_vsdinv _19305_ (.A(\cpuregs[2][16] ),
    .Y(_00778_));
 sky130_vsdinv _19306_ (.A(\cpuregs[3][16] ),
    .Y(_00779_));
 sky130_vsdinv _19307_ (.A(\cpuregs[4][16] ),
    .Y(_00781_));
 sky130_vsdinv _19308_ (.A(\cpuregs[5][16] ),
    .Y(_00782_));
 sky130_vsdinv _19309_ (.A(\cpuregs[6][16] ),
    .Y(_00783_));
 sky130_vsdinv _19310_ (.A(\cpuregs[7][16] ),
    .Y(_00784_));
 sky130_vsdinv _19311_ (.A(\cpuregs[8][16] ),
    .Y(_00786_));
 sky130_vsdinv _19312_ (.A(\cpuregs[9][16] ),
    .Y(_00787_));
 sky130_vsdinv _19313_ (.A(\cpuregs[10][16] ),
    .Y(_00788_));
 sky130_vsdinv _19314_ (.A(\cpuregs[11][16] ),
    .Y(_00789_));
 sky130_vsdinv _19315_ (.A(\cpuregs[12][16] ),
    .Y(_00791_));
 sky130_vsdinv _19316_ (.A(\cpuregs[13][16] ),
    .Y(_00792_));
 sky130_vsdinv _19317_ (.A(\cpuregs[14][16] ),
    .Y(_00793_));
 sky130_vsdinv _19318_ (.A(\cpuregs[15][16] ),
    .Y(_00794_));
 sky130_vsdinv _19319_ (.A(\cpuregs[16][16] ),
    .Y(_00797_));
 sky130_vsdinv _19320_ (.A(\cpuregs[17][16] ),
    .Y(_00798_));
 sky130_vsdinv _19321_ (.A(\cpuregs[18][16] ),
    .Y(_00799_));
 sky130_vsdinv _19322_ (.A(\cpuregs[19][16] ),
    .Y(_00800_));
 sky130_vsdinv _19323_ (.A(\cpuregs[0][17] ),
    .Y(_00803_));
 sky130_vsdinv _19324_ (.A(\cpuregs[1][17] ),
    .Y(_00804_));
 sky130_vsdinv _19325_ (.A(\cpuregs[2][17] ),
    .Y(_00805_));
 sky130_vsdinv _19326_ (.A(\cpuregs[3][17] ),
    .Y(_00806_));
 sky130_vsdinv _19327_ (.A(\cpuregs[4][17] ),
    .Y(_00808_));
 sky130_vsdinv _19328_ (.A(\cpuregs[5][17] ),
    .Y(_00809_));
 sky130_vsdinv _19329_ (.A(\cpuregs[6][17] ),
    .Y(_00810_));
 sky130_vsdinv _19330_ (.A(\cpuregs[7][17] ),
    .Y(_00811_));
 sky130_vsdinv _19331_ (.A(\cpuregs[8][17] ),
    .Y(_00813_));
 sky130_vsdinv _19332_ (.A(\cpuregs[9][17] ),
    .Y(_00814_));
 sky130_vsdinv _19333_ (.A(\cpuregs[10][17] ),
    .Y(_00815_));
 sky130_vsdinv _19334_ (.A(\cpuregs[11][17] ),
    .Y(_00816_));
 sky130_vsdinv _19335_ (.A(\cpuregs[12][17] ),
    .Y(_00818_));
 sky130_vsdinv _19336_ (.A(\cpuregs[13][17] ),
    .Y(_00819_));
 sky130_vsdinv _19337_ (.A(\cpuregs[14][17] ),
    .Y(_00820_));
 sky130_vsdinv _19338_ (.A(\cpuregs[15][17] ),
    .Y(_00821_));
 sky130_vsdinv _19339_ (.A(\cpuregs[16][17] ),
    .Y(_00824_));
 sky130_vsdinv _19340_ (.A(\cpuregs[17][17] ),
    .Y(_00825_));
 sky130_vsdinv _19341_ (.A(\cpuregs[18][17] ),
    .Y(_00826_));
 sky130_vsdinv _19342_ (.A(\cpuregs[19][17] ),
    .Y(_00827_));
 sky130_vsdinv _19343_ (.A(\cpuregs[0][18] ),
    .Y(_00830_));
 sky130_vsdinv _19344_ (.A(\cpuregs[1][18] ),
    .Y(_00831_));
 sky130_vsdinv _19345_ (.A(\cpuregs[2][18] ),
    .Y(_00832_));
 sky130_vsdinv _19346_ (.A(\cpuregs[3][18] ),
    .Y(_00833_));
 sky130_vsdinv _19347_ (.A(\cpuregs[4][18] ),
    .Y(_00835_));
 sky130_vsdinv _19348_ (.A(\cpuregs[5][18] ),
    .Y(_00836_));
 sky130_vsdinv _19349_ (.A(\cpuregs[6][18] ),
    .Y(_00837_));
 sky130_vsdinv _19350_ (.A(\cpuregs[7][18] ),
    .Y(_00838_));
 sky130_vsdinv _19351_ (.A(\cpuregs[8][18] ),
    .Y(_00840_));
 sky130_vsdinv _19352_ (.A(\cpuregs[9][18] ),
    .Y(_00841_));
 sky130_vsdinv _19353_ (.A(\cpuregs[10][18] ),
    .Y(_00842_));
 sky130_vsdinv _19354_ (.A(\cpuregs[11][18] ),
    .Y(_00843_));
 sky130_vsdinv _19355_ (.A(\cpuregs[12][18] ),
    .Y(_00845_));
 sky130_vsdinv _19356_ (.A(\cpuregs[13][18] ),
    .Y(_00846_));
 sky130_vsdinv _19357_ (.A(\cpuregs[14][18] ),
    .Y(_00847_));
 sky130_vsdinv _19358_ (.A(\cpuregs[15][18] ),
    .Y(_00848_));
 sky130_vsdinv _19359_ (.A(\cpuregs[16][18] ),
    .Y(_00851_));
 sky130_vsdinv _19360_ (.A(\cpuregs[17][18] ),
    .Y(_00852_));
 sky130_vsdinv _19361_ (.A(\cpuregs[18][18] ),
    .Y(_00853_));
 sky130_vsdinv _19362_ (.A(\cpuregs[19][18] ),
    .Y(_00854_));
 sky130_vsdinv _19363_ (.A(\cpuregs[0][19] ),
    .Y(_00857_));
 sky130_vsdinv _19364_ (.A(\cpuregs[1][19] ),
    .Y(_00858_));
 sky130_vsdinv _19365_ (.A(\cpuregs[2][19] ),
    .Y(_00859_));
 sky130_vsdinv _19366_ (.A(\cpuregs[3][19] ),
    .Y(_00860_));
 sky130_vsdinv _19367_ (.A(\cpuregs[4][19] ),
    .Y(_00862_));
 sky130_vsdinv _19368_ (.A(\cpuregs[5][19] ),
    .Y(_00863_));
 sky130_vsdinv _19369_ (.A(\cpuregs[6][19] ),
    .Y(_00864_));
 sky130_vsdinv _19370_ (.A(\cpuregs[7][19] ),
    .Y(_00865_));
 sky130_vsdinv _19371_ (.A(\cpuregs[8][19] ),
    .Y(_00867_));
 sky130_vsdinv _19372_ (.A(\cpuregs[9][19] ),
    .Y(_00868_));
 sky130_vsdinv _19373_ (.A(\cpuregs[10][19] ),
    .Y(_00869_));
 sky130_vsdinv _19374_ (.A(\cpuregs[11][19] ),
    .Y(_00870_));
 sky130_vsdinv _19375_ (.A(\cpuregs[12][19] ),
    .Y(_00872_));
 sky130_vsdinv _19376_ (.A(\cpuregs[13][19] ),
    .Y(_00873_));
 sky130_vsdinv _19377_ (.A(\cpuregs[14][19] ),
    .Y(_00874_));
 sky130_vsdinv _19378_ (.A(\cpuregs[15][19] ),
    .Y(_00875_));
 sky130_vsdinv _19379_ (.A(\cpuregs[16][19] ),
    .Y(_00878_));
 sky130_vsdinv _19380_ (.A(\cpuregs[17][19] ),
    .Y(_00879_));
 sky130_vsdinv _19381_ (.A(\cpuregs[18][19] ),
    .Y(_00880_));
 sky130_vsdinv _19382_ (.A(\cpuregs[19][19] ),
    .Y(_00881_));
 sky130_vsdinv _19383_ (.A(\cpuregs[0][20] ),
    .Y(_00884_));
 sky130_vsdinv _19384_ (.A(\cpuregs[1][20] ),
    .Y(_00885_));
 sky130_vsdinv _19385_ (.A(\cpuregs[2][20] ),
    .Y(_00886_));
 sky130_vsdinv _19386_ (.A(\cpuregs[3][20] ),
    .Y(_00887_));
 sky130_vsdinv _19387_ (.A(\cpuregs[4][20] ),
    .Y(_00889_));
 sky130_vsdinv _19388_ (.A(\cpuregs[5][20] ),
    .Y(_00890_));
 sky130_vsdinv _19389_ (.A(\cpuregs[6][20] ),
    .Y(_00891_));
 sky130_vsdinv _19390_ (.A(\cpuregs[7][20] ),
    .Y(_00892_));
 sky130_vsdinv _19391_ (.A(\cpuregs[8][20] ),
    .Y(_00894_));
 sky130_vsdinv _19392_ (.A(\cpuregs[9][20] ),
    .Y(_00895_));
 sky130_vsdinv _19393_ (.A(\cpuregs[10][20] ),
    .Y(_00896_));
 sky130_vsdinv _19394_ (.A(\cpuregs[11][20] ),
    .Y(_00897_));
 sky130_vsdinv _19395_ (.A(\cpuregs[12][20] ),
    .Y(_00899_));
 sky130_vsdinv _19396_ (.A(\cpuregs[13][20] ),
    .Y(_00900_));
 sky130_vsdinv _19397_ (.A(\cpuregs[14][20] ),
    .Y(_00901_));
 sky130_vsdinv _19398_ (.A(\cpuregs[15][20] ),
    .Y(_00902_));
 sky130_vsdinv _19399_ (.A(\cpuregs[16][20] ),
    .Y(_00905_));
 sky130_vsdinv _19400_ (.A(\cpuregs[17][20] ),
    .Y(_00906_));
 sky130_vsdinv _19401_ (.A(\cpuregs[18][20] ),
    .Y(_00907_));
 sky130_vsdinv _19402_ (.A(\cpuregs[19][20] ),
    .Y(_00908_));
 sky130_vsdinv _19403_ (.A(\cpuregs[0][21] ),
    .Y(_00911_));
 sky130_vsdinv _19404_ (.A(\cpuregs[1][21] ),
    .Y(_00912_));
 sky130_vsdinv _19405_ (.A(\cpuregs[2][21] ),
    .Y(_00913_));
 sky130_vsdinv _19406_ (.A(\cpuregs[3][21] ),
    .Y(_00914_));
 sky130_vsdinv _19407_ (.A(\cpuregs[4][21] ),
    .Y(_00916_));
 sky130_vsdinv _19408_ (.A(\cpuregs[5][21] ),
    .Y(_00917_));
 sky130_vsdinv _19409_ (.A(\cpuregs[6][21] ),
    .Y(_00918_));
 sky130_vsdinv _19410_ (.A(\cpuregs[7][21] ),
    .Y(_00919_));
 sky130_fd_sc_hd__clkbuf_4 _19411_ (.A(_14264_),
    .X(_14828_));
 sky130_fd_sc_hd__clkbuf_4 _19412_ (.A(_14268_),
    .X(_14829_));
 sky130_fd_sc_hd__nor2_8 _19413_ (.A(_14828_),
    .B(_14829_),
    .Y(_00304_));
 sky130_vsdinv _19414_ (.A(\cpuregs[8][21] ),
    .Y(_00921_));
 sky130_vsdinv _19415_ (.A(\cpuregs[9][21] ),
    .Y(_00922_));
 sky130_vsdinv _19416_ (.A(\cpuregs[10][21] ),
    .Y(_00923_));
 sky130_vsdinv _19417_ (.A(\cpuregs[11][21] ),
    .Y(_00924_));
 sky130_vsdinv _19418_ (.A(\cpuregs[12][21] ),
    .Y(_00926_));
 sky130_vsdinv _19419_ (.A(\cpuregs[13][21] ),
    .Y(_00927_));
 sky130_vsdinv _19420_ (.A(\cpuregs[14][21] ),
    .Y(_00928_));
 sky130_vsdinv _19421_ (.A(\cpuregs[15][21] ),
    .Y(_00929_));
 sky130_vsdinv _19422_ (.A(\cpuregs[16][21] ),
    .Y(_00932_));
 sky130_vsdinv _19423_ (.A(\cpuregs[17][21] ),
    .Y(_00933_));
 sky130_vsdinv _19424_ (.A(\cpuregs[18][21] ),
    .Y(_00934_));
 sky130_vsdinv _19425_ (.A(\cpuregs[19][21] ),
    .Y(_00935_));
 sky130_vsdinv _19426_ (.A(\cpuregs[0][22] ),
    .Y(_00938_));
 sky130_vsdinv _19427_ (.A(\cpuregs[1][22] ),
    .Y(_00939_));
 sky130_vsdinv _19428_ (.A(\cpuregs[2][22] ),
    .Y(_00940_));
 sky130_vsdinv _19429_ (.A(\cpuregs[3][22] ),
    .Y(_00941_));
 sky130_vsdinv _19430_ (.A(\cpuregs[4][22] ),
    .Y(_00943_));
 sky130_vsdinv _19431_ (.A(\cpuregs[5][22] ),
    .Y(_00944_));
 sky130_vsdinv _19432_ (.A(\cpuregs[6][22] ),
    .Y(_00945_));
 sky130_vsdinv _19433_ (.A(\cpuregs[7][22] ),
    .Y(_00946_));
 sky130_fd_sc_hd__and4_1 _19434_ (.A(_14696_),
    .B(_12648_),
    .C(instr_lw),
    .D(_12651_),
    .X(_14830_));
 sky130_fd_sc_hd__a21oi_1 _19435_ (.A1(instr_sw),
    .A2(_14814_),
    .B1(_14830_),
    .Y(_14831_));
 sky130_fd_sc_hd__or2b_1 _19436_ (.A(_14821_),
    .B_N(\mem_wordsize[0] ),
    .X(_14832_));
 sky130_fd_sc_hd__o221ai_1 _19437_ (.A1(_12964_),
    .A2(_00322_),
    .B1(_00296_),
    .B2(_14831_),
    .C1(_14832_),
    .Y(_00045_));
 sky130_vsdinv _19438_ (.A(\cpuregs[8][22] ),
    .Y(_00948_));
 sky130_vsdinv _19439_ (.A(\cpuregs[9][22] ),
    .Y(_00949_));
 sky130_vsdinv _19440_ (.A(\cpuregs[10][22] ),
    .Y(_00950_));
 sky130_vsdinv _19441_ (.A(\cpuregs[11][22] ),
    .Y(_00951_));
 sky130_vsdinv _19442_ (.A(\cpuregs[12][22] ),
    .Y(_00953_));
 sky130_vsdinv _19443_ (.A(\cpuregs[13][22] ),
    .Y(_00954_));
 sky130_vsdinv _19444_ (.A(\cpuregs[14][22] ),
    .Y(_00955_));
 sky130_vsdinv _19445_ (.A(\cpuregs[15][22] ),
    .Y(_00956_));
 sky130_vsdinv _19446_ (.A(\cpuregs[16][22] ),
    .Y(_00959_));
 sky130_vsdinv _19447_ (.A(\cpuregs[17][22] ),
    .Y(_00960_));
 sky130_vsdinv _19448_ (.A(\cpuregs[18][22] ),
    .Y(_00961_));
 sky130_vsdinv _19449_ (.A(\cpuregs[19][22] ),
    .Y(_00962_));
 sky130_vsdinv _19450_ (.A(\cpuregs[0][23] ),
    .Y(_00965_));
 sky130_vsdinv _19451_ (.A(\cpuregs[1][23] ),
    .Y(_00966_));
 sky130_vsdinv _19452_ (.A(\cpuregs[2][23] ),
    .Y(_00967_));
 sky130_vsdinv _19453_ (.A(\cpuregs[3][23] ),
    .Y(_00968_));
 sky130_vsdinv _19454_ (.A(\cpuregs[4][23] ),
    .Y(_00970_));
 sky130_vsdinv _19455_ (.A(\cpuregs[5][23] ),
    .Y(_00971_));
 sky130_vsdinv _19456_ (.A(\cpuregs[6][23] ),
    .Y(_00972_));
 sky130_vsdinv _19457_ (.A(\cpuregs[7][23] ),
    .Y(_00973_));
 sky130_vsdinv _19458_ (.A(\cpuregs[8][23] ),
    .Y(_00975_));
 sky130_vsdinv _19459_ (.A(\cpuregs[9][23] ),
    .Y(_00976_));
 sky130_vsdinv _19460_ (.A(\cpuregs[10][23] ),
    .Y(_00977_));
 sky130_vsdinv _19461_ (.A(\cpuregs[11][23] ),
    .Y(_00978_));
 sky130_vsdinv _19462_ (.A(\cpuregs[12][23] ),
    .Y(_00980_));
 sky130_vsdinv _19463_ (.A(\cpuregs[13][23] ),
    .Y(_00981_));
 sky130_vsdinv _19464_ (.A(\cpuregs[14][23] ),
    .Y(_00982_));
 sky130_vsdinv _19465_ (.A(\cpuregs[15][23] ),
    .Y(_00983_));
 sky130_vsdinv _19466_ (.A(\cpuregs[16][23] ),
    .Y(_00986_));
 sky130_vsdinv _19467_ (.A(\cpuregs[17][23] ),
    .Y(_00987_));
 sky130_vsdinv _19468_ (.A(\cpuregs[18][23] ),
    .Y(_00988_));
 sky130_vsdinv _19469_ (.A(\cpuregs[19][23] ),
    .Y(_00989_));
 sky130_vsdinv _19470_ (.A(\cpuregs[0][24] ),
    .Y(_00992_));
 sky130_vsdinv _19471_ (.A(\cpuregs[1][24] ),
    .Y(_00993_));
 sky130_vsdinv _19472_ (.A(\cpuregs[2][24] ),
    .Y(_00994_));
 sky130_vsdinv _19473_ (.A(\cpuregs[3][24] ),
    .Y(_00995_));
 sky130_vsdinv _19474_ (.A(\cpuregs[4][24] ),
    .Y(_00997_));
 sky130_vsdinv _19475_ (.A(\cpuregs[5][24] ),
    .Y(_00998_));
 sky130_vsdinv _19476_ (.A(\cpuregs[6][24] ),
    .Y(_00999_));
 sky130_vsdinv _19477_ (.A(\cpuregs[7][24] ),
    .Y(_01000_));
 sky130_vsdinv _19478_ (.A(\cpuregs[8][24] ),
    .Y(_01002_));
 sky130_vsdinv _19479_ (.A(\cpuregs[9][24] ),
    .Y(_01003_));
 sky130_vsdinv _19480_ (.A(\cpuregs[10][24] ),
    .Y(_01004_));
 sky130_vsdinv _19481_ (.A(\cpuregs[11][24] ),
    .Y(_01005_));
 sky130_vsdinv _19482_ (.A(\cpuregs[12][24] ),
    .Y(_01007_));
 sky130_vsdinv _19483_ (.A(\cpuregs[13][24] ),
    .Y(_01008_));
 sky130_vsdinv _19484_ (.A(\cpuregs[14][24] ),
    .Y(_01009_));
 sky130_vsdinv _19485_ (.A(\cpuregs[15][24] ),
    .Y(_01010_));
 sky130_vsdinv _19486_ (.A(\cpuregs[16][24] ),
    .Y(_01013_));
 sky130_vsdinv _19487_ (.A(\cpuregs[17][24] ),
    .Y(_01014_));
 sky130_vsdinv _19488_ (.A(\cpuregs[18][24] ),
    .Y(_01015_));
 sky130_vsdinv _19489_ (.A(\cpuregs[19][24] ),
    .Y(_01016_));
 sky130_vsdinv _19490_ (.A(\cpuregs[0][25] ),
    .Y(_01019_));
 sky130_vsdinv _19491_ (.A(\cpuregs[1][25] ),
    .Y(_01020_));
 sky130_vsdinv _19492_ (.A(\cpuregs[2][25] ),
    .Y(_01021_));
 sky130_vsdinv _19493_ (.A(\cpuregs[3][25] ),
    .Y(_01022_));
 sky130_vsdinv _19494_ (.A(\cpuregs[4][25] ),
    .Y(_01024_));
 sky130_vsdinv _19495_ (.A(\cpuregs[5][25] ),
    .Y(_01025_));
 sky130_vsdinv _19496_ (.A(\cpuregs[6][25] ),
    .Y(_01026_));
 sky130_vsdinv _19497_ (.A(\cpuregs[7][25] ),
    .Y(_01027_));
 sky130_fd_sc_hd__nor2b_1 _19498_ (.A(\mem_state[1] ),
    .B_N(_12631_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _19499_ (.A(_12676_),
    .B(_00289_),
    .Y(_00298_));
 sky130_vsdinv _19500_ (.A(\cpuregs[8][25] ),
    .Y(_01029_));
 sky130_vsdinv _19501_ (.A(\cpuregs[9][25] ),
    .Y(_01030_));
 sky130_vsdinv _19502_ (.A(\cpuregs[10][25] ),
    .Y(_01031_));
 sky130_vsdinv _19503_ (.A(\cpuregs[11][25] ),
    .Y(_01032_));
 sky130_vsdinv _19504_ (.A(\cpuregs[12][25] ),
    .Y(_01034_));
 sky130_vsdinv _19505_ (.A(\cpuregs[13][25] ),
    .Y(_01035_));
 sky130_vsdinv _19506_ (.A(\cpuregs[14][25] ),
    .Y(_01036_));
 sky130_vsdinv _19507_ (.A(\cpuregs[15][25] ),
    .Y(_01037_));
 sky130_vsdinv _19508_ (.A(\cpuregs[16][25] ),
    .Y(_01040_));
 sky130_vsdinv _19509_ (.A(\cpuregs[17][25] ),
    .Y(_01041_));
 sky130_vsdinv _19510_ (.A(\cpuregs[18][25] ),
    .Y(_01042_));
 sky130_vsdinv _19511_ (.A(\cpuregs[19][25] ),
    .Y(_01043_));
 sky130_vsdinv _19512_ (.A(\cpuregs[0][26] ),
    .Y(_01046_));
 sky130_vsdinv _19513_ (.A(\cpuregs[1][26] ),
    .Y(_01047_));
 sky130_vsdinv _19514_ (.A(\cpuregs[2][26] ),
    .Y(_01048_));
 sky130_vsdinv _19515_ (.A(\cpuregs[3][26] ),
    .Y(_01049_));
 sky130_vsdinv _19516_ (.A(\cpuregs[4][26] ),
    .Y(_01051_));
 sky130_vsdinv _19517_ (.A(\cpuregs[5][26] ),
    .Y(_01052_));
 sky130_vsdinv _19518_ (.A(\cpuregs[6][26] ),
    .Y(_01053_));
 sky130_vsdinv _19519_ (.A(\cpuregs[7][26] ),
    .Y(_01054_));
 sky130_vsdinv _19520_ (.A(\cpuregs[8][26] ),
    .Y(_01056_));
 sky130_vsdinv _19521_ (.A(\cpuregs[9][26] ),
    .Y(_01057_));
 sky130_vsdinv _19522_ (.A(\cpuregs[10][26] ),
    .Y(_01058_));
 sky130_vsdinv _19523_ (.A(\cpuregs[11][26] ),
    .Y(_01059_));
 sky130_vsdinv _19524_ (.A(\cpuregs[12][26] ),
    .Y(_01061_));
 sky130_vsdinv _19525_ (.A(\cpuregs[13][26] ),
    .Y(_01062_));
 sky130_vsdinv _19526_ (.A(\cpuregs[14][26] ),
    .Y(_01063_));
 sky130_vsdinv _19527_ (.A(\cpuregs[15][26] ),
    .Y(_01064_));
 sky130_vsdinv _19528_ (.A(\cpuregs[16][26] ),
    .Y(_01067_));
 sky130_vsdinv _19529_ (.A(\cpuregs[17][26] ),
    .Y(_01068_));
 sky130_vsdinv _19530_ (.A(\cpuregs[18][26] ),
    .Y(_01069_));
 sky130_vsdinv _19531_ (.A(\cpuregs[19][26] ),
    .Y(_01070_));
 sky130_fd_sc_hd__inv_2 _19532_ (.A(\mem_wordsize[1] ),
    .Y(_14833_));
 sky130_fd_sc_hd__and3b_1 _19533_ (.A_N(_12976_),
    .B(instr_sb),
    .C(_14212_),
    .X(_14834_));
 sky130_fd_sc_hd__o211a_1 _19534_ (.A1(instr_lbu),
    .A2(instr_lb),
    .B1(_12651_),
    .C1(_14696_),
    .X(_14835_));
 sky130_fd_sc_hd__o21a_1 _19535_ (.A1(_14834_),
    .A2(_14835_),
    .B1(_12644_),
    .X(_14836_));
 sky130_fd_sc_hd__o21bai_1 _19536_ (.A1(_14833_),
    .A2(_14821_),
    .B1_N(_14836_),
    .Y(_00046_));
 sky130_vsdinv _19537_ (.A(\cpuregs[0][27] ),
    .Y(_01073_));
 sky130_vsdinv _19538_ (.A(\cpuregs[1][27] ),
    .Y(_01074_));
 sky130_vsdinv _19539_ (.A(\cpuregs[2][27] ),
    .Y(_01075_));
 sky130_vsdinv _19540_ (.A(\cpuregs[3][27] ),
    .Y(_01076_));
 sky130_vsdinv _19541_ (.A(\cpuregs[4][27] ),
    .Y(_01078_));
 sky130_vsdinv _19542_ (.A(\cpuregs[5][27] ),
    .Y(_01079_));
 sky130_vsdinv _19543_ (.A(\cpuregs[6][27] ),
    .Y(_01080_));
 sky130_vsdinv _19544_ (.A(\cpuregs[7][27] ),
    .Y(_01081_));
 sky130_vsdinv _19545_ (.A(\cpuregs[8][27] ),
    .Y(_01083_));
 sky130_vsdinv _19546_ (.A(\cpuregs[9][27] ),
    .Y(_01084_));
 sky130_vsdinv _19547_ (.A(\cpuregs[10][27] ),
    .Y(_01085_));
 sky130_vsdinv _19548_ (.A(\cpuregs[11][27] ),
    .Y(_01086_));
 sky130_vsdinv _19549_ (.A(\cpuregs[12][27] ),
    .Y(_01088_));
 sky130_vsdinv _19550_ (.A(\cpuregs[13][27] ),
    .Y(_01089_));
 sky130_vsdinv _19551_ (.A(\cpuregs[14][27] ),
    .Y(_01090_));
 sky130_vsdinv _19552_ (.A(\cpuregs[15][27] ),
    .Y(_01091_));
 sky130_vsdinv _19553_ (.A(\cpuregs[16][27] ),
    .Y(_01094_));
 sky130_vsdinv _19554_ (.A(\cpuregs[17][27] ),
    .Y(_01095_));
 sky130_vsdinv _19555_ (.A(\cpuregs[18][27] ),
    .Y(_01096_));
 sky130_vsdinv _19556_ (.A(\cpuregs[19][27] ),
    .Y(_01097_));
 sky130_vsdinv _19557_ (.A(\cpuregs[0][28] ),
    .Y(_01100_));
 sky130_vsdinv _19558_ (.A(\cpuregs[1][28] ),
    .Y(_01101_));
 sky130_vsdinv _19559_ (.A(\cpuregs[2][28] ),
    .Y(_01102_));
 sky130_vsdinv _19560_ (.A(\cpuregs[3][28] ),
    .Y(_01103_));
 sky130_vsdinv _19561_ (.A(\cpuregs[4][28] ),
    .Y(_01105_));
 sky130_vsdinv _19562_ (.A(\cpuregs[5][28] ),
    .Y(_01106_));
 sky130_vsdinv _19563_ (.A(\cpuregs[6][28] ),
    .Y(_01107_));
 sky130_vsdinv _19564_ (.A(\cpuregs[7][28] ),
    .Y(_01108_));
 sky130_vsdinv _19565_ (.A(\cpuregs[8][28] ),
    .Y(_01110_));
 sky130_vsdinv _19566_ (.A(\cpuregs[9][28] ),
    .Y(_01111_));
 sky130_vsdinv _19567_ (.A(\cpuregs[10][28] ),
    .Y(_01112_));
 sky130_vsdinv _19568_ (.A(\cpuregs[11][28] ),
    .Y(_01113_));
 sky130_vsdinv _19569_ (.A(\cpuregs[12][28] ),
    .Y(_01115_));
 sky130_vsdinv _19570_ (.A(\cpuregs[13][28] ),
    .Y(_01116_));
 sky130_vsdinv _19571_ (.A(\cpuregs[14][28] ),
    .Y(_01117_));
 sky130_vsdinv _19572_ (.A(\cpuregs[15][28] ),
    .Y(_01118_));
 sky130_vsdinv _19573_ (.A(\cpuregs[16][28] ),
    .Y(_01121_));
 sky130_vsdinv _19574_ (.A(\cpuregs[17][28] ),
    .Y(_01122_));
 sky130_vsdinv _19575_ (.A(\cpuregs[18][28] ),
    .Y(_01123_));
 sky130_vsdinv _19576_ (.A(\cpuregs[19][28] ),
    .Y(_01124_));
 sky130_vsdinv _19577_ (.A(\cpuregs[0][29] ),
    .Y(_01127_));
 sky130_vsdinv _19578_ (.A(\cpuregs[1][29] ),
    .Y(_01128_));
 sky130_vsdinv _19579_ (.A(\cpuregs[2][29] ),
    .Y(_01129_));
 sky130_vsdinv _19580_ (.A(\cpuregs[3][29] ),
    .Y(_01130_));
 sky130_vsdinv _19581_ (.A(\cpuregs[4][29] ),
    .Y(_01132_));
 sky130_vsdinv _19582_ (.A(\cpuregs[5][29] ),
    .Y(_01133_));
 sky130_vsdinv _19583_ (.A(\cpuregs[6][29] ),
    .Y(_01134_));
 sky130_vsdinv _19584_ (.A(\cpuregs[7][29] ),
    .Y(_01135_));
 sky130_vsdinv _19585_ (.A(\cpuregs[8][29] ),
    .Y(_01137_));
 sky130_vsdinv _19586_ (.A(\cpuregs[9][29] ),
    .Y(_01138_));
 sky130_vsdinv _19587_ (.A(\cpuregs[10][29] ),
    .Y(_01139_));
 sky130_vsdinv _19588_ (.A(\cpuregs[11][29] ),
    .Y(_01140_));
 sky130_vsdinv _19589_ (.A(\cpuregs[12][29] ),
    .Y(_01142_));
 sky130_vsdinv _19590_ (.A(\cpuregs[13][29] ),
    .Y(_01143_));
 sky130_fd_sc_hd__clkbuf_4 _19591_ (.A(_14536_),
    .X(_14837_));
 sky130_fd_sc_hd__and2_1 _19592_ (.A(_14837_),
    .B(_00294_),
    .X(_00295_));
 sky130_vsdinv _19593_ (.A(\cpuregs[14][29] ),
    .Y(_01144_));
 sky130_vsdinv _19594_ (.A(\cpuregs[15][29] ),
    .Y(_01145_));
 sky130_vsdinv _19595_ (.A(\cpuregs[16][29] ),
    .Y(_01148_));
 sky130_vsdinv _19596_ (.A(\cpuregs[17][29] ),
    .Y(_01149_));
 sky130_vsdinv _19597_ (.A(\cpuregs[18][29] ),
    .Y(_01150_));
 sky130_vsdinv _19598_ (.A(\cpuregs[19][29] ),
    .Y(_01151_));
 sky130_vsdinv _19599_ (.A(\cpuregs[0][30] ),
    .Y(_01154_));
 sky130_vsdinv _19600_ (.A(\cpuregs[1][30] ),
    .Y(_01155_));
 sky130_vsdinv _19601_ (.A(\cpuregs[2][30] ),
    .Y(_01156_));
 sky130_vsdinv _19602_ (.A(\cpuregs[3][30] ),
    .Y(_01157_));
 sky130_vsdinv _19603_ (.A(\cpuregs[4][30] ),
    .Y(_01159_));
 sky130_vsdinv _19604_ (.A(\cpuregs[5][30] ),
    .Y(_01160_));
 sky130_vsdinv _19605_ (.A(\cpuregs[6][30] ),
    .Y(_01161_));
 sky130_vsdinv _19606_ (.A(\cpuregs[7][30] ),
    .Y(_01162_));
 sky130_vsdinv _19607_ (.A(\cpuregs[8][30] ),
    .Y(_01164_));
 sky130_vsdinv _19608_ (.A(\cpuregs[9][30] ),
    .Y(_01165_));
 sky130_vsdinv _19609_ (.A(\cpuregs[10][30] ),
    .Y(_01166_));
 sky130_vsdinv _19610_ (.A(\cpuregs[11][30] ),
    .Y(_01167_));
 sky130_vsdinv _19611_ (.A(\cpuregs[12][30] ),
    .Y(_01169_));
 sky130_vsdinv _19612_ (.A(\cpuregs[13][30] ),
    .Y(_01170_));
 sky130_vsdinv _19613_ (.A(\cpuregs[14][30] ),
    .Y(_01171_));
 sky130_vsdinv _19614_ (.A(\cpuregs[15][30] ),
    .Y(_01172_));
 sky130_vsdinv _19615_ (.A(\cpuregs[16][30] ),
    .Y(_01175_));
 sky130_vsdinv _19616_ (.A(\cpuregs[17][30] ),
    .Y(_01176_));
 sky130_vsdinv _19617_ (.A(\cpuregs[18][30] ),
    .Y(_01177_));
 sky130_vsdinv _19618_ (.A(\cpuregs[19][30] ),
    .Y(_01178_));
 sky130_vsdinv _19619_ (.A(\cpuregs[0][31] ),
    .Y(_01181_));
 sky130_vsdinv _19620_ (.A(\cpuregs[1][31] ),
    .Y(_01182_));
 sky130_vsdinv _19621_ (.A(\cpuregs[2][31] ),
    .Y(_01183_));
 sky130_vsdinv _19622_ (.A(\cpuregs[3][31] ),
    .Y(_01184_));
 sky130_vsdinv _19623_ (.A(\cpuregs[4][31] ),
    .Y(_01186_));
 sky130_vsdinv _19624_ (.A(\cpuregs[5][31] ),
    .Y(_01187_));
 sky130_vsdinv _19625_ (.A(\cpuregs[6][31] ),
    .Y(_01188_));
 sky130_vsdinv _19626_ (.A(\cpuregs[7][31] ),
    .Y(_01189_));
 sky130_vsdinv _19627_ (.A(\cpuregs[8][31] ),
    .Y(_01191_));
 sky130_vsdinv _19628_ (.A(\cpuregs[9][31] ),
    .Y(_01192_));
 sky130_vsdinv _19629_ (.A(\cpuregs[10][31] ),
    .Y(_01193_));
 sky130_vsdinv _19630_ (.A(\cpuregs[11][31] ),
    .Y(_01194_));
 sky130_vsdinv _19631_ (.A(\cpuregs[12][31] ),
    .Y(_01196_));
 sky130_vsdinv _19632_ (.A(\cpuregs[13][31] ),
    .Y(_01197_));
 sky130_vsdinv _19633_ (.A(\cpuregs[14][31] ),
    .Y(_01198_));
 sky130_vsdinv _19634_ (.A(\cpuregs[15][31] ),
    .Y(_01199_));
 sky130_vsdinv _19635_ (.A(\cpuregs[16][31] ),
    .Y(_01202_));
 sky130_vsdinv _19636_ (.A(\cpuregs[17][31] ),
    .Y(_01203_));
 sky130_vsdinv _19637_ (.A(\cpuregs[18][31] ),
    .Y(_01204_));
 sky130_vsdinv _19638_ (.A(\cpuregs[19][31] ),
    .Y(_01205_));
 sky130_fd_sc_hd__or2_4 _19639_ (.A(\timer[27] ),
    .B(\timer[26] ),
    .X(_14838_));
 sky130_fd_sc_hd__nor2_4 _19640_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .Y(_14839_));
 sky130_vsdinv _19641_ (.A(\timer[31] ),
    .Y(_14840_));
 sky130_fd_sc_hd__nand3b_4 _19642_ (.A_N(\timer[30] ),
    .B(_14839_),
    .C(_14840_),
    .Y(_14841_));
 sky130_fd_sc_hd__or4_4 _19643_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(\timer[23] ),
    .D(\timer[22] ),
    .X(_14842_));
 sky130_fd_sc_hd__or2_4 _19644_ (.A(\timer[25] ),
    .B(\timer[24] ),
    .X(_14843_));
 sky130_fd_sc_hd__or2_4 _19645_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .X(_14844_));
 sky130_fd_sc_hd__nor2_4 _19646_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .Y(_14845_));
 sky130_vsdinv _19647_ (.A(\timer[3] ),
    .Y(_14846_));
 sky130_vsdinv _19648_ (.A(\timer[2] ),
    .Y(_14847_));
 sky130_fd_sc_hd__nand3_4 _19649_ (.A(_14845_),
    .B(_14846_),
    .C(_14847_),
    .Y(_14848_));
 sky130_fd_sc_hd__nor3_4 _19650_ (.A(\timer[6] ),
    .B(_14844_),
    .C(_14848_),
    .Y(_14849_));
 sky130_vsdinv _19651_ (.A(\timer[7] ),
    .Y(_14850_));
 sky130_fd_sc_hd__nor3_1 _19652_ (.A(\timer[9] ),
    .B(\timer[8] ),
    .C(\timer[11] ),
    .Y(_14851_));
 sky130_fd_sc_hd__and2b_1 _19653_ (.A_N(\timer[10] ),
    .B(_14851_),
    .X(_14852_));
 sky130_fd_sc_hd__nand3_2 _19654_ (.A(_14849_),
    .B(_14850_),
    .C(_14852_),
    .Y(_14853_));
 sky130_fd_sc_hd__nor2_1 _19655_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .Y(_14854_));
 sky130_fd_sc_hd__nor3b_4 _19656_ (.A(\timer[15] ),
    .B(\timer[14] ),
    .C_N(_14854_),
    .Y(_14855_));
 sky130_fd_sc_hd__or2_4 _19657_ (.A(\timer[17] ),
    .B(\timer[16] ),
    .X(_14856_));
 sky130_fd_sc_hd__nor3_4 _19658_ (.A(\timer[19] ),
    .B(\timer[18] ),
    .C(_14856_),
    .Y(_14857_));
 sky130_fd_sc_hd__nand3b_4 _19659_ (.A_N(_14853_),
    .B(_14855_),
    .C(_14857_),
    .Y(_14858_));
 sky130_fd_sc_hd__nor3_4 _19660_ (.A(_14842_),
    .B(_14843_),
    .C(_14858_),
    .Y(_14859_));
 sky130_fd_sc_hd__nor3b_4 _19661_ (.A(_14838_),
    .B(_14841_),
    .C_N(_14859_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _19662_ (.A(\timer[0] ),
    .B(net417),
    .Y(_01209_));
 sky130_fd_sc_hd__xnor2_1 _19663_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .Y(_01211_));
 sky130_fd_sc_hd__xor2_1 _19664_ (.A(\timer[2] ),
    .B(_14845_),
    .X(_01214_));
 sky130_fd_sc_hd__nor3_4 _19665_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .C(\timer[2] ),
    .Y(_14860_));
 sky130_fd_sc_hd__xor2_1 _19666_ (.A(\timer[3] ),
    .B(_14860_),
    .X(_01217_));
 sky130_vsdinv _19667_ (.A(\timer[4] ),
    .Y(_14861_));
 sky130_fd_sc_hd__xor2_1 _19668_ (.A(_14861_),
    .B(_14848_),
    .X(_01220_));
 sky130_fd_sc_hd__nand3_1 _19669_ (.A(_14860_),
    .B(_14846_),
    .C(_14861_),
    .Y(_14862_));
 sky130_fd_sc_hd__o2bb2ai_1 _19670_ (.A1_N(\timer[5] ),
    .A2_N(_14862_),
    .B1(_14844_),
    .B2(_14848_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor2_4 _19671_ (.A(_14844_),
    .B(_14848_),
    .Y(_14863_));
 sky130_fd_sc_hd__xor2_1 _19672_ (.A(\timer[6] ),
    .B(_14863_),
    .X(_01226_));
 sky130_fd_sc_hd__xor2_1 _19673_ (.A(\timer[7] ),
    .B(_14849_),
    .X(_01229_));
 sky130_fd_sc_hd__nand3b_4 _19674_ (.A_N(\timer[6] ),
    .B(_14863_),
    .C(_14850_),
    .Y(_14864_));
 sky130_fd_sc_hd__xnor2_1 _19675_ (.A(\timer[8] ),
    .B(_14864_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand3b_4 _19676_ (.A_N(\timer[8] ),
    .B(_14849_),
    .C(_14850_),
    .Y(_14865_));
 sky130_fd_sc_hd__xnor2_1 _19677_ (.A(\timer[9] ),
    .B(_14865_),
    .Y(_01235_));
 sky130_fd_sc_hd__nor3_2 _19678_ (.A(\timer[9] ),
    .B(\timer[8] ),
    .C(_14864_),
    .Y(_14866_));
 sky130_fd_sc_hd__xor2_1 _19679_ (.A(\timer[10] ),
    .B(_14866_),
    .X(_01238_));
 sky130_fd_sc_hd__nor3_2 _19680_ (.A(\timer[9] ),
    .B(\timer[10] ),
    .C(_14865_),
    .Y(_14867_));
 sky130_fd_sc_hd__xor2_1 _19681_ (.A(\timer[11] ),
    .B(_14867_),
    .X(_01241_));
 sky130_fd_sc_hd__buf_4 _19682_ (.A(_14853_),
    .X(_14868_));
 sky130_fd_sc_hd__xnor2_1 _19683_ (.A(\timer[12] ),
    .B(_14868_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _19684_ (.A(\timer[12] ),
    .B(_14868_),
    .Y(_14869_));
 sky130_fd_sc_hd__xor2_1 _19685_ (.A(\timer[13] ),
    .B(_14869_),
    .X(_01247_));
 sky130_fd_sc_hd__nor3_2 _19686_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .C(_14868_),
    .Y(_14870_));
 sky130_fd_sc_hd__xor2_1 _19687_ (.A(\timer[14] ),
    .B(_14870_),
    .X(_01250_));
 sky130_fd_sc_hd__nor3b_4 _19688_ (.A(\timer[14] ),
    .B(_14868_),
    .C_N(_14854_),
    .Y(_14871_));
 sky130_fd_sc_hd__xor2_1 _19689_ (.A(\timer[15] ),
    .B(_14871_),
    .X(_01253_));
 sky130_fd_sc_hd__and4_2 _19690_ (.A(_14849_),
    .B(_14850_),
    .C(_14852_),
    .D(_14855_),
    .X(_14872_));
 sky130_fd_sc_hd__xor2_1 _19691_ (.A(\timer[16] ),
    .B(_14872_),
    .X(_01256_));
 sky130_fd_sc_hd__nor3b_4 _19692_ (.A(\timer[16] ),
    .B(_14868_),
    .C_N(_14855_),
    .Y(_14873_));
 sky130_fd_sc_hd__xor2_1 _19693_ (.A(\timer[17] ),
    .B(_14873_),
    .X(_01259_));
 sky130_fd_sc_hd__nor3b_4 _19694_ (.A(_14856_),
    .B(_14868_),
    .C_N(_14855_),
    .Y(_14874_));
 sky130_fd_sc_hd__xor2_1 _19695_ (.A(\timer[18] ),
    .B(_14874_),
    .X(_01262_));
 sky130_fd_sc_hd__nor3b_4 _19696_ (.A(\timer[18] ),
    .B(_14856_),
    .C_N(_14872_),
    .Y(_14875_));
 sky130_fd_sc_hd__xor2_1 _19697_ (.A(\timer[19] ),
    .B(_14875_),
    .X(_01265_));
 sky130_fd_sc_hd__xnor2_1 _19698_ (.A(\timer[20] ),
    .B(_14858_),
    .Y(_01268_));
 sky130_fd_sc_hd__nand3b_4 _19699_ (.A_N(\timer[20] ),
    .B(_14872_),
    .C(_14857_),
    .Y(_14876_));
 sky130_fd_sc_hd__xnor2_1 _19700_ (.A(\timer[21] ),
    .B(_14876_),
    .Y(_01271_));
 sky130_fd_sc_hd__nor3_4 _19701_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(_14858_),
    .Y(_14877_));
 sky130_fd_sc_hd__xor2_1 _19702_ (.A(\timer[22] ),
    .B(_14877_),
    .X(_01274_));
 sky130_fd_sc_hd__nor3_4 _19703_ (.A(\timer[21] ),
    .B(\timer[22] ),
    .C(_14876_),
    .Y(_14878_));
 sky130_fd_sc_hd__xor2_1 _19704_ (.A(\timer[23] ),
    .B(_14878_),
    .X(_01277_));
 sky130_fd_sc_hd__nor2_2 _19705_ (.A(_14842_),
    .B(_14858_),
    .Y(_14879_));
 sky130_fd_sc_hd__xor2_1 _19706_ (.A(\timer[24] ),
    .B(_14879_),
    .X(_01280_));
 sky130_fd_sc_hd__nor3_4 _19707_ (.A(\timer[24] ),
    .B(_14842_),
    .C(_14858_),
    .Y(_14880_));
 sky130_fd_sc_hd__xor2_1 _19708_ (.A(\timer[25] ),
    .B(_14880_),
    .X(_01283_));
 sky130_fd_sc_hd__xor2_1 _19709_ (.A(\timer[26] ),
    .B(_14859_),
    .X(_01286_));
 sky130_fd_sc_hd__nor3b_4 _19710_ (.A(\timer[26] ),
    .B(_14843_),
    .C_N(_14879_),
    .Y(_14881_));
 sky130_fd_sc_hd__xor2_1 _19711_ (.A(\timer[27] ),
    .B(_14881_),
    .X(_01289_));
 sky130_fd_sc_hd__nor3b_4 _19712_ (.A(_14843_),
    .B(_14838_),
    .C_N(_14879_),
    .Y(_14882_));
 sky130_fd_sc_hd__xor2_1 _19713_ (.A(\timer[28] ),
    .B(_14882_),
    .X(_01292_));
 sky130_fd_sc_hd__nor3b_4 _19714_ (.A(\timer[28] ),
    .B(_14838_),
    .C_N(_14859_),
    .Y(_14883_));
 sky130_fd_sc_hd__xor2_1 _19715_ (.A(\timer[29] ),
    .B(_14883_),
    .X(_01295_));
 sky130_fd_sc_hd__nor3b_4 _19716_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .C_N(_14882_),
    .Y(_14884_));
 sky130_fd_sc_hd__xor2_1 _19717_ (.A(\timer[30] ),
    .B(_14884_),
    .X(_01298_));
 sky130_fd_sc_hd__nand3b_2 _19718_ (.A_N(\timer[30] ),
    .B(_14882_),
    .C(_14839_),
    .Y(_14885_));
 sky130_fd_sc_hd__xor2_1 _19719_ (.A(_14840_),
    .B(_14885_),
    .X(_01301_));
 sky130_fd_sc_hd__clkbuf_2 _19720_ (.A(_14121_),
    .X(_14886_));
 sky130_fd_sc_hd__nor2b_1 _19721_ (.A(_14886_),
    .B_N(\decoded_imm[5] ),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2b_1 _19722_ (.A(_14886_),
    .B_N(_14563_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2b_1 _19723_ (.A(_14886_),
    .B_N(_14566_),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2b_1 _19724_ (.A(_14886_),
    .B_N(_14569_),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2b_1 _19725_ (.A(_14886_),
    .B_N(_14571_),
    .Y(_01323_));
 sky130_fd_sc_hd__nor2b_1 _19726_ (.A(_14886_),
    .B_N(\decoded_imm[10] ),
    .Y(_01325_));
 sky130_fd_sc_hd__clkbuf_2 _19727_ (.A(_14121_),
    .X(_14887_));
 sky130_fd_sc_hd__nor2b_1 _19728_ (.A(_14887_),
    .B_N(\decoded_imm[11] ),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2b_1 _19729_ (.A(_14887_),
    .B_N(\decoded_imm[12] ),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2b_1 _19730_ (.A(_14887_),
    .B_N(\decoded_imm[13] ),
    .Y(_01331_));
 sky130_fd_sc_hd__nor2b_1 _19731_ (.A(_14887_),
    .B_N(\decoded_imm[14] ),
    .Y(_01333_));
 sky130_fd_sc_hd__nor2b_1 _19732_ (.A(_14887_),
    .B_N(\decoded_imm[15] ),
    .Y(_01335_));
 sky130_fd_sc_hd__nor2b_1 _19733_ (.A(_14887_),
    .B_N(_14594_),
    .Y(_01337_));
 sky130_fd_sc_hd__buf_2 _19734_ (.A(is_slli_srli_srai),
    .X(_14888_));
 sky130_fd_sc_hd__nor2b_1 _19735_ (.A(_14888_),
    .B_N(_14597_),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2b_1 _19736_ (.A(_14888_),
    .B_N(_14600_),
    .Y(_01341_));
 sky130_fd_sc_hd__nor2b_1 _19737_ (.A(_14888_),
    .B_N(\decoded_imm[19] ),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2b_1 _19738_ (.A(_14888_),
    .B_N(\decoded_imm[20] ),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2b_1 _19739_ (.A(_14888_),
    .B_N(\decoded_imm[21] ),
    .Y(_01347_));
 sky130_fd_sc_hd__nor2b_1 _19740_ (.A(_14888_),
    .B_N(\decoded_imm[22] ),
    .Y(_01349_));
 sky130_fd_sc_hd__clkbuf_2 _19741_ (.A(is_slli_srli_srai),
    .X(_14889_));
 sky130_fd_sc_hd__nor2b_1 _19742_ (.A(_14889_),
    .B_N(\decoded_imm[23] ),
    .Y(_01351_));
 sky130_fd_sc_hd__nor2b_1 _19743_ (.A(_14889_),
    .B_N(_14615_),
    .Y(_01353_));
 sky130_fd_sc_hd__nor2b_1 _19744_ (.A(_14889_),
    .B_N(_14618_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2b_1 _19745_ (.A(_14889_),
    .B_N(_14620_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2b_1 _19746_ (.A(_14889_),
    .B_N(_14623_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2b_1 _19747_ (.A(_14889_),
    .B_N(_14625_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2b_1 _19748_ (.A(_14121_),
    .B_N(\decoded_imm[29] ),
    .Y(_01363_));
 sky130_fd_sc_hd__nor2b_1 _19749_ (.A(_14121_),
    .B_N(\decoded_imm[30] ),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2b_1 _19750_ (.A(_14121_),
    .B_N(\decoded_imm[31] ),
    .Y(_01367_));
 sky130_fd_sc_hd__buf_2 _19751_ (.A(_14205_),
    .X(_14890_));
 sky130_fd_sc_hd__nor2b_1 _19752_ (.A(_14890_),
    .B_N(\reg_next_pc[0] ),
    .Y(_01369_));
 sky130_fd_sc_hd__xor2_1 _19753_ (.A(\decoded_imm[0] ),
    .B(_14269_),
    .X(_01371_));
 sky130_fd_sc_hd__nor2b_1 _19754_ (.A(_14890_),
    .B_N(\reg_pc[1] ),
    .Y(_01372_));
 sky130_fd_sc_hd__and2_1 _19755_ (.A(\decoded_imm[0] ),
    .B(_14268_),
    .X(_14891_));
 sky130_fd_sc_hd__xnor2_2 _19756_ (.A(net317),
    .B(\decoded_imm[1] ),
    .Y(_14892_));
 sky130_fd_sc_hd__xnor2_1 _19757_ (.A(_14891_),
    .B(_14892_),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2b_1 _19758_ (.A(_14890_),
    .B_N(_13249_),
    .Y(_01375_));
 sky130_fd_sc_hd__xor2_1 _19759_ (.A(_14262_),
    .B(\decoded_imm[2] ),
    .X(_14893_));
 sky130_fd_sc_hd__nand3b_4 _19760_ (.A_N(_14892_),
    .B(\decoded_imm[0] ),
    .C(net306),
    .Y(_14894_));
 sky130_fd_sc_hd__nand2_1 _19761_ (.A(net317),
    .B(\decoded_imm[1] ),
    .Y(_14895_));
 sky130_fd_sc_hd__nand2_1 _19762_ (.A(_14894_),
    .B(_14895_),
    .Y(_14896_));
 sky130_fd_sc_hd__xor2_1 _19763_ (.A(_14893_),
    .B(_14896_),
    .X(_01377_));
 sky130_fd_sc_hd__nor2b_1 _19764_ (.A(_14890_),
    .B_N(_13246_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_1 _19765_ (.A(net331),
    .B(\decoded_imm[3] ),
    .Y(_14897_));
 sky130_fd_sc_hd__and2_1 _19766_ (.A(net331),
    .B(\decoded_imm[3] ),
    .X(_14898_));
 sky130_fd_sc_hd__nor2_1 _19767_ (.A(_14897_),
    .B(_14898_),
    .Y(_14899_));
 sky130_fd_sc_hd__o2bb2ai_1 _19768_ (.A1_N(_14895_),
    .A2_N(_14894_),
    .B1(_14261_),
    .B2(\decoded_imm[2] ),
    .Y(_14900_));
 sky130_fd_sc_hd__nand2_1 _19769_ (.A(_14261_),
    .B(\decoded_imm[2] ),
    .Y(_14901_));
 sky130_fd_sc_hd__nand2_1 _19770_ (.A(_14900_),
    .B(_14901_),
    .Y(_14902_));
 sky130_fd_sc_hd__xor2_1 _19771_ (.A(_14899_),
    .B(_14902_),
    .X(_01380_));
 sky130_fd_sc_hd__nor2b_1 _19772_ (.A(_14890_),
    .B_N(_13244_),
    .Y(_01381_));
 sky130_fd_sc_hd__xor2_1 _19773_ (.A(_14259_),
    .B(\decoded_imm[4] ),
    .X(_14903_));
 sky130_vsdinv _19774_ (.A(_14897_),
    .Y(_14904_));
 sky130_fd_sc_hd__a21o_1 _19775_ (.A1(_14902_),
    .A2(_14904_),
    .B1(_14898_),
    .X(_14905_));
 sky130_fd_sc_hd__xor2_1 _19776_ (.A(_14903_),
    .B(_14905_),
    .X(_01383_));
 sky130_fd_sc_hd__nor2b_1 _19777_ (.A(_14890_),
    .B_N(_13241_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_1 _19778_ (.A(net333),
    .B(\decoded_imm[5] ),
    .Y(_14906_));
 sky130_fd_sc_hd__and2_1 _19779_ (.A(net333),
    .B(\decoded_imm[5] ),
    .X(_14907_));
 sky130_fd_sc_hd__nor2_1 _19780_ (.A(_14906_),
    .B(_14907_),
    .Y(_14908_));
 sky130_fd_sc_hd__o21ai_1 _19781_ (.A1(_14258_),
    .A2(\decoded_imm[4] ),
    .B1(_14905_),
    .Y(_14909_));
 sky130_fd_sc_hd__nand2_1 _19782_ (.A(_14258_),
    .B(\decoded_imm[4] ),
    .Y(_14910_));
 sky130_fd_sc_hd__nand2_1 _19783_ (.A(_14909_),
    .B(_14910_),
    .Y(_14911_));
 sky130_fd_sc_hd__xor2_1 _19784_ (.A(_14908_),
    .B(_14911_),
    .X(_01386_));
 sky130_fd_sc_hd__clkbuf_2 _19785_ (.A(_14205_),
    .X(_14912_));
 sky130_fd_sc_hd__nor2b_1 _19786_ (.A(_14912_),
    .B_N(_13237_),
    .Y(_01387_));
 sky130_fd_sc_hd__xor2_4 _19787_ (.A(_14255_),
    .B(_14563_),
    .X(_14913_));
 sky130_vsdinv _19788_ (.A(_14906_),
    .Y(_14914_));
 sky130_fd_sc_hd__a21o_1 _19789_ (.A1(_14911_),
    .A2(_14914_),
    .B1(_14907_),
    .X(_14915_));
 sky130_fd_sc_hd__xor2_1 _19790_ (.A(_14913_),
    .B(_14915_),
    .X(_01389_));
 sky130_fd_sc_hd__nor2b_1 _19791_ (.A(_14912_),
    .B_N(\reg_pc[7] ),
    .Y(_01390_));
 sky130_fd_sc_hd__xnor2_1 _19792_ (.A(net335),
    .B(\decoded_imm[7] ),
    .Y(_14916_));
 sky130_fd_sc_hd__and2_1 _19793_ (.A(_14256_),
    .B(_14563_),
    .X(_14917_));
 sky130_fd_sc_hd__a21oi_1 _19794_ (.A1(_14915_),
    .A2(_14913_),
    .B1(_14917_),
    .Y(_14918_));
 sky130_fd_sc_hd__xor2_1 _19795_ (.A(_14916_),
    .B(_14918_),
    .X(_01392_));
 sky130_fd_sc_hd__nor2b_1 _19796_ (.A(_14912_),
    .B_N(\reg_pc[8] ),
    .Y(_01393_));
 sky130_fd_sc_hd__xor2_2 _19797_ (.A(_14250_),
    .B(\decoded_imm[8] ),
    .X(_14919_));
 sky130_fd_sc_hd__and2b_1 _19798_ (.A_N(_14916_),
    .B(_14913_),
    .X(_14920_));
 sky130_fd_sc_hd__o211a_1 _19799_ (.A1(_14252_),
    .A2(_14566_),
    .B1(_14255_),
    .C1(_14563_),
    .X(_14921_));
 sky130_fd_sc_hd__a221oi_2 _19800_ (.A1(_14252_),
    .A2(_14566_),
    .B1(_14915_),
    .B2(_14920_),
    .C1(_14921_),
    .Y(_14922_));
 sky130_fd_sc_hd__xnor2_1 _19801_ (.A(_14919_),
    .B(_14922_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor2b_1 _19802_ (.A(_14912_),
    .B_N(_13229_),
    .Y(_01396_));
 sky130_fd_sc_hd__xnor2_2 _19803_ (.A(_14248_),
    .B(\decoded_imm[9] ),
    .Y(_14923_));
 sky130_fd_sc_hd__and2b_1 _19804_ (.A_N(_14922_),
    .B(_14919_),
    .X(_14924_));
 sky130_fd_sc_hd__a21oi_1 _19805_ (.A1(_14251_),
    .A2(_14569_),
    .B1(_14924_),
    .Y(_14925_));
 sky130_fd_sc_hd__xor2_1 _19806_ (.A(_14923_),
    .B(_14925_),
    .X(_01398_));
 sky130_fd_sc_hd__nor2b_1 _19807_ (.A(_14912_),
    .B_N(_13226_),
    .Y(_01399_));
 sky130_fd_sc_hd__xor2_2 _19808_ (.A(net307),
    .B(\decoded_imm[10] ),
    .X(_14926_));
 sky130_fd_sc_hd__o211a_1 _19809_ (.A1(_14248_),
    .A2(_14571_),
    .B1(_14250_),
    .C1(_14569_),
    .X(_14927_));
 sky130_fd_sc_hd__nor3b_2 _19810_ (.A(_14923_),
    .B(_14922_),
    .C_N(_14919_),
    .Y(_14928_));
 sky130_fd_sc_hd__a211o_1 _19811_ (.A1(_14248_),
    .A2(_14571_),
    .B1(_14927_),
    .C1(_14928_),
    .X(_14929_));
 sky130_fd_sc_hd__xor2_1 _19812_ (.A(_14926_),
    .B(_14929_),
    .X(_01401_));
 sky130_fd_sc_hd__nor2b_1 _19813_ (.A(_14912_),
    .B_N(_13223_),
    .Y(_01402_));
 sky130_fd_sc_hd__xor2_2 _19814_ (.A(net308),
    .B(\decoded_imm[11] ),
    .X(_14930_));
 sky130_fd_sc_hd__and2_1 _19815_ (.A(net307),
    .B(\decoded_imm[10] ),
    .X(_14931_));
 sky130_fd_sc_hd__a21o_1 _19816_ (.A1(_14929_),
    .A2(_14926_),
    .B1(_14931_),
    .X(_14932_));
 sky130_fd_sc_hd__xor2_1 _19817_ (.A(_14930_),
    .B(_14932_),
    .X(_01404_));
 sky130_fd_sc_hd__clkbuf_2 _19818_ (.A(_14205_),
    .X(_14933_));
 sky130_fd_sc_hd__nor2b_1 _19819_ (.A(_14933_),
    .B_N(\reg_pc[12] ),
    .Y(_01405_));
 sky130_fd_sc_hd__xor2_2 _19820_ (.A(net309),
    .B(\decoded_imm[12] ),
    .X(_14934_));
 sky130_fd_sc_hd__and2_1 _19821_ (.A(net308),
    .B(\decoded_imm[11] ),
    .X(_14935_));
 sky130_fd_sc_hd__a21o_1 _19822_ (.A1(_14932_),
    .A2(_14930_),
    .B1(_14935_),
    .X(_14936_));
 sky130_fd_sc_hd__xor2_1 _19823_ (.A(_14934_),
    .B(_14936_),
    .X(_01407_));
 sky130_fd_sc_hd__nor2b_1 _19824_ (.A(_14933_),
    .B_N(_13215_),
    .Y(_01408_));
 sky130_fd_sc_hd__xor2_2 _19825_ (.A(net310),
    .B(\decoded_imm[13] ),
    .X(_14937_));
 sky130_fd_sc_hd__and2_1 _19826_ (.A(net309),
    .B(\decoded_imm[12] ),
    .X(_14938_));
 sky130_fd_sc_hd__a21o_1 _19827_ (.A1(_14936_),
    .A2(_14934_),
    .B1(_14938_),
    .X(_14939_));
 sky130_fd_sc_hd__xor2_1 _19828_ (.A(_14937_),
    .B(_14939_),
    .X(_01410_));
 sky130_fd_sc_hd__nor2b_1 _19829_ (.A(_14933_),
    .B_N(_13213_),
    .Y(_01411_));
 sky130_fd_sc_hd__xor2_2 _19830_ (.A(net311),
    .B(\decoded_imm[14] ),
    .X(_14940_));
 sky130_fd_sc_hd__and2_1 _19831_ (.A(net310),
    .B(\decoded_imm[13] ),
    .X(_14941_));
 sky130_fd_sc_hd__a21o_1 _19832_ (.A1(_14939_),
    .A2(_14937_),
    .B1(_14941_),
    .X(_14942_));
 sky130_fd_sc_hd__xor2_1 _19833_ (.A(_14940_),
    .B(_14942_),
    .X(_01413_));
 sky130_fd_sc_hd__nor2b_1 _19834_ (.A(_14933_),
    .B_N(_13208_),
    .Y(_01414_));
 sky130_fd_sc_hd__xnor2_2 _19835_ (.A(net312),
    .B(\decoded_imm[15] ),
    .Y(_14943_));
 sky130_fd_sc_hd__and2_1 _19836_ (.A(net311),
    .B(\decoded_imm[14] ),
    .X(_14944_));
 sky130_fd_sc_hd__a21oi_2 _19837_ (.A1(_14942_),
    .A2(_14940_),
    .B1(_14944_),
    .Y(_14945_));
 sky130_fd_sc_hd__xor2_1 _19838_ (.A(_14943_),
    .B(_14945_),
    .X(_01416_));
 sky130_fd_sc_hd__nor2b_1 _19839_ (.A(_14933_),
    .B_N(_13205_),
    .Y(_01417_));
 sky130_fd_sc_hd__xor2_4 _19840_ (.A(net313),
    .B(\decoded_imm[16] ),
    .X(_14946_));
 sky130_fd_sc_hd__and2_1 _19841_ (.A(net312),
    .B(\decoded_imm[15] ),
    .X(_14947_));
 sky130_fd_sc_hd__o21bai_2 _19842_ (.A1(_14943_),
    .A2(_14945_),
    .B1_N(_14947_),
    .Y(_14948_));
 sky130_fd_sc_hd__xor2_1 _19843_ (.A(_14946_),
    .B(_14948_),
    .X(_01419_));
 sky130_fd_sc_hd__nor2b_1 _19844_ (.A(_14933_),
    .B_N(_13203_),
    .Y(_01420_));
 sky130_fd_sc_hd__xnor2_1 _19845_ (.A(net314),
    .B(_14597_),
    .Y(_14949_));
 sky130_fd_sc_hd__and2_1 _19846_ (.A(_14240_),
    .B(_14594_),
    .X(_14950_));
 sky130_fd_sc_hd__a21oi_1 _19847_ (.A1(_14948_),
    .A2(_14946_),
    .B1(_14950_),
    .Y(_14951_));
 sky130_fd_sc_hd__xor2_1 _19848_ (.A(_14949_),
    .B(_14951_),
    .X(_01422_));
 sky130_fd_sc_hd__buf_2 _19849_ (.A(instr_lui),
    .X(_14952_));
 sky130_fd_sc_hd__nor2b_1 _19850_ (.A(_14952_),
    .B_N(_13199_),
    .Y(_01423_));
 sky130_fd_sc_hd__xnor2_1 _19851_ (.A(net315),
    .B(_14600_),
    .Y(_14953_));
 sky130_fd_sc_hd__and2b_1 _19852_ (.A_N(_14949_),
    .B(_14946_),
    .X(_14954_));
 sky130_fd_sc_hd__o211a_1 _19853_ (.A1(_14237_),
    .A2(_14597_),
    .B1(_14239_),
    .C1(_14594_),
    .X(_14955_));
 sky130_fd_sc_hd__a221oi_2 _19854_ (.A1(_14237_),
    .A2(_14597_),
    .B1(_14948_),
    .B2(_14954_),
    .C1(_14955_),
    .Y(_14956_));
 sky130_fd_sc_hd__xor2_1 _19855_ (.A(_14953_),
    .B(_14956_),
    .X(_01425_));
 sky130_fd_sc_hd__nor2b_1 _19856_ (.A(_14952_),
    .B_N(_13194_),
    .Y(_01426_));
 sky130_fd_sc_hd__xor2_4 _19857_ (.A(net316),
    .B(\decoded_imm[19] ),
    .X(_14957_));
 sky130_fd_sc_hd__and2_1 _19858_ (.A(net315),
    .B(_14600_),
    .X(_14958_));
 sky130_fd_sc_hd__o21bai_2 _19859_ (.A1(_14953_),
    .A2(_14956_),
    .B1_N(_14958_),
    .Y(_14959_));
 sky130_fd_sc_hd__xor2_1 _19860_ (.A(_14957_),
    .B(_14959_),
    .X(_01428_));
 sky130_fd_sc_hd__nor2b_1 _19861_ (.A(_14952_),
    .B_N(_13192_),
    .Y(_01429_));
 sky130_fd_sc_hd__xnor2_1 _19862_ (.A(net318),
    .B(\decoded_imm[20] ),
    .Y(_14960_));
 sky130_fd_sc_hd__and2_1 _19863_ (.A(net316),
    .B(\decoded_imm[19] ),
    .X(_14961_));
 sky130_fd_sc_hd__a21oi_4 _19864_ (.A1(_14959_),
    .A2(_14957_),
    .B1(_14961_),
    .Y(_14962_));
 sky130_fd_sc_hd__xor2_1 _19865_ (.A(_14960_),
    .B(_14962_),
    .X(_01431_));
 sky130_fd_sc_hd__nor2b_1 _19866_ (.A(_14952_),
    .B_N(_13189_),
    .Y(_01432_));
 sky130_fd_sc_hd__xor2_2 _19867_ (.A(net319),
    .B(\decoded_imm[21] ),
    .X(_14963_));
 sky130_fd_sc_hd__and2_1 _19868_ (.A(net318),
    .B(\decoded_imm[20] ),
    .X(_14964_));
 sky130_fd_sc_hd__o21bai_2 _19869_ (.A1(_14960_),
    .A2(_14962_),
    .B1_N(_14964_),
    .Y(_14965_));
 sky130_fd_sc_hd__xor2_1 _19870_ (.A(_14963_),
    .B(_14965_),
    .X(_01434_));
 sky130_fd_sc_hd__nor2b_1 _19871_ (.A(_14952_),
    .B_N(_13186_),
    .Y(_01435_));
 sky130_fd_sc_hd__xnor2_1 _19872_ (.A(net320),
    .B(\decoded_imm[22] ),
    .Y(_14966_));
 sky130_fd_sc_hd__and2_1 _19873_ (.A(net319),
    .B(\decoded_imm[21] ),
    .X(_14967_));
 sky130_fd_sc_hd__a21oi_2 _19874_ (.A1(_14965_),
    .A2(_14963_),
    .B1(_14967_),
    .Y(_14968_));
 sky130_fd_sc_hd__xor2_1 _19875_ (.A(_14966_),
    .B(_14968_),
    .X(_01437_));
 sky130_fd_sc_hd__nor2b_1 _19876_ (.A(_14952_),
    .B_N(_13182_),
    .Y(_01438_));
 sky130_fd_sc_hd__xor2_4 _19877_ (.A(net321),
    .B(\decoded_imm[23] ),
    .X(_14969_));
 sky130_fd_sc_hd__and2_1 _19878_ (.A(net320),
    .B(\decoded_imm[22] ),
    .X(_14970_));
 sky130_fd_sc_hd__o21bai_2 _19879_ (.A1(_14966_),
    .A2(_14968_),
    .B1_N(_14970_),
    .Y(_14971_));
 sky130_fd_sc_hd__xor2_1 _19880_ (.A(_14969_),
    .B(_14971_),
    .X(_01440_));
 sky130_fd_sc_hd__clkbuf_2 _19881_ (.A(instr_lui),
    .X(_14972_));
 sky130_fd_sc_hd__nor2b_1 _19882_ (.A(_14972_),
    .B_N(\reg_pc[24] ),
    .Y(_01441_));
 sky130_fd_sc_hd__xor2_4 _19883_ (.A(_14228_),
    .B(_14615_),
    .X(_14973_));
 sky130_fd_sc_hd__and2_1 _19884_ (.A(net321),
    .B(\decoded_imm[23] ),
    .X(_14974_));
 sky130_fd_sc_hd__a21oi_4 _19885_ (.A1(_14971_),
    .A2(_14969_),
    .B1(_14974_),
    .Y(_14975_));
 sky130_fd_sc_hd__xnor2_1 _19886_ (.A(_14973_),
    .B(_14975_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2b_1 _19887_ (.A(_14972_),
    .B_N(_13175_),
    .Y(_01444_));
 sky130_fd_sc_hd__xor2_2 _19888_ (.A(_14225_),
    .B(_14618_),
    .X(_14976_));
 sky130_fd_sc_hd__and2b_1 _19889_ (.A_N(_14975_),
    .B(_14973_),
    .X(_14977_));
 sky130_fd_sc_hd__a21oi_1 _19890_ (.A1(_14229_),
    .A2(_14615_),
    .B1(_14977_),
    .Y(_14978_));
 sky130_fd_sc_hd__xnor2_1 _19891_ (.A(_14976_),
    .B(_14978_),
    .Y(_01446_));
 sky130_fd_sc_hd__nor2b_1 _19892_ (.A(_14972_),
    .B_N(_13173_),
    .Y(_01447_));
 sky130_fd_sc_hd__xor2_2 _19893_ (.A(_14223_),
    .B(\decoded_imm[26] ),
    .X(_14979_));
 sky130_fd_sc_hd__nand2_1 _19894_ (.A(_14973_),
    .B(_14976_),
    .Y(_14980_));
 sky130_fd_sc_hd__and2_1 _19895_ (.A(_14225_),
    .B(_14618_),
    .X(_14981_));
 sky130_vsdinv _19896_ (.A(_14981_),
    .Y(_14982_));
 sky130_fd_sc_hd__o211ai_2 _19897_ (.A1(_14226_),
    .A2(_14618_),
    .B1(_14228_),
    .C1(_14615_),
    .Y(_14983_));
 sky130_fd_sc_hd__o211ai_4 _19898_ (.A1(_14980_),
    .A2(_14975_),
    .B1(_14982_),
    .C1(_14983_),
    .Y(_14984_));
 sky130_fd_sc_hd__xor2_1 _19899_ (.A(_14979_),
    .B(_14984_),
    .X(_01449_));
 sky130_fd_sc_hd__nor2b_1 _19900_ (.A(_14972_),
    .B_N(_13170_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_1 _19901_ (.A(_14221_),
    .B(_14623_),
    .Y(_14985_));
 sky130_fd_sc_hd__and2_1 _19902_ (.A(_14221_),
    .B(\decoded_imm[27] ),
    .X(_14986_));
 sky130_fd_sc_hd__nor2_1 _19903_ (.A(_14985_),
    .B(_14986_),
    .Y(_14987_));
 sky130_fd_sc_hd__and2_1 _19904_ (.A(_14224_),
    .B(_14620_),
    .X(_14988_));
 sky130_fd_sc_hd__a21oi_1 _19905_ (.A1(_14984_),
    .A2(_14979_),
    .B1(_14988_),
    .Y(_14989_));
 sky130_fd_sc_hd__xnor2_1 _19906_ (.A(_14987_),
    .B(_14989_),
    .Y(_01452_));
 sky130_fd_sc_hd__nor2b_1 _19907_ (.A(_14972_),
    .B_N(\reg_pc[28] ),
    .Y(_01453_));
 sky130_fd_sc_hd__xnor2_1 _19908_ (.A(_14220_),
    .B(_14625_),
    .Y(_14990_));
 sky130_fd_sc_hd__and2_1 _19909_ (.A(_14979_),
    .B(_14987_),
    .X(_14991_));
 sky130_fd_sc_hd__o211a_1 _19910_ (.A1(_14222_),
    .A2(_14623_),
    .B1(_14223_),
    .C1(_14620_),
    .X(_14992_));
 sky130_fd_sc_hd__nor2_1 _19911_ (.A(_14986_),
    .B(_14992_),
    .Y(_14993_));
 sky130_fd_sc_hd__a21boi_4 _19912_ (.A1(_14984_),
    .A2(_14991_),
    .B1_N(_14993_),
    .Y(_14994_));
 sky130_fd_sc_hd__xor2_1 _19913_ (.A(_14990_),
    .B(_14994_),
    .X(_01455_));
 sky130_fd_sc_hd__nor2b_1 _19914_ (.A(_14972_),
    .B_N(_13159_),
    .Y(_01456_));
 sky130_fd_sc_hd__xor2_1 _19915_ (.A(_14218_),
    .B(\decoded_imm[29] ),
    .X(_14995_));
 sky130_fd_sc_hd__nor2_1 _19916_ (.A(_14219_),
    .B(_14625_),
    .Y(_14996_));
 sky130_fd_sc_hd__and2_1 _19917_ (.A(_14219_),
    .B(_14625_),
    .X(_14997_));
 sky130_fd_sc_hd__o21bai_2 _19918_ (.A1(_14996_),
    .A2(_14994_),
    .B1_N(_14997_),
    .Y(_14998_));
 sky130_fd_sc_hd__xor2_1 _19919_ (.A(_14995_),
    .B(_14998_),
    .X(_01458_));
 sky130_fd_sc_hd__nor2b_1 _19920_ (.A(_14205_),
    .B_N(\reg_pc[30] ),
    .Y(_01459_));
 sky130_fd_sc_hd__xnor2_2 _19921_ (.A(net329),
    .B(\decoded_imm[30] ),
    .Y(_14999_));
 sky130_vsdinv _19922_ (.A(net327),
    .Y(_15000_));
 sky130_fd_sc_hd__nand2_1 _19923_ (.A(_15000_),
    .B(_14627_),
    .Y(_15001_));
 sky130_fd_sc_hd__and2_1 _19924_ (.A(_14218_),
    .B(\decoded_imm[29] ),
    .X(_15002_));
 sky130_fd_sc_hd__a21oi_4 _19925_ (.A1(_14998_),
    .A2(_15001_),
    .B1(_15002_),
    .Y(_15003_));
 sky130_fd_sc_hd__xor2_1 _19926_ (.A(_14999_),
    .B(_15003_),
    .X(_01461_));
 sky130_fd_sc_hd__nor2b_1 _19927_ (.A(_14205_),
    .B_N(\reg_pc[31] ),
    .Y(_01462_));
 sky130_fd_sc_hd__and2_1 _19928_ (.A(_14217_),
    .B(\decoded_imm[30] ),
    .X(_15004_));
 sky130_fd_sc_hd__nor2_1 _19929_ (.A(_14999_),
    .B(_15003_),
    .Y(_15005_));
 sky130_fd_sc_hd__xnor2_1 _19930_ (.A(net330),
    .B(\decoded_imm[31] ),
    .Y(_15006_));
 sky130_vsdinv _19931_ (.A(_15006_),
    .Y(_15007_));
 sky130_fd_sc_hd__o21bai_1 _19932_ (.A1(_15004_),
    .A2(_15005_),
    .B1_N(_15007_),
    .Y(_15008_));
 sky130_vsdinv _19933_ (.A(_15004_),
    .Y(_15009_));
 sky130_fd_sc_hd__o211ai_1 _19934_ (.A1(_14999_),
    .A2(_15003_),
    .B1(_15009_),
    .C1(_15007_),
    .Y(_15010_));
 sky130_fd_sc_hd__nand2_1 _19935_ (.A(_15008_),
    .B(_15010_),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_1 _19936_ (.A(_14837_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__and2_1 _19937_ (.A(_14837_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__inv_2 _19938_ (.A(\reg_next_pc[4] ),
    .Y(_01471_));
 sky130_fd_sc_hd__buf_2 _19939_ (.A(_12878_),
    .X(_15011_));
 sky130_fd_sc_hd__a21oi_1 _19940_ (.A1(_14837_),
    .A2(_01473_),
    .B1(_15011_),
    .Y(_01474_));
 sky130_fd_sc_hd__and2_1 _19941_ (.A(_14837_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__clkbuf_2 _19942_ (.A(_14536_),
    .X(_15012_));
 sky130_fd_sc_hd__and2_1 _19943_ (.A(_15012_),
    .B(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__and2_1 _19944_ (.A(_15012_),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__and2_1 _19945_ (.A(_15012_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__and2_1 _19946_ (.A(_15012_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__and2_1 _19947_ (.A(_15012_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__and2_1 _19948_ (.A(_15012_),
    .B(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__clkbuf_2 _19949_ (.A(_12663_),
    .X(_15013_));
 sky130_fd_sc_hd__and2_1 _19950_ (.A(_15013_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__and2_1 _19951_ (.A(_15013_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__and2_1 _19952_ (.A(_15013_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__and2_1 _19953_ (.A(_15013_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__and2_1 _19954_ (.A(_15013_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__and2_1 _19955_ (.A(_15013_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__buf_1 _19956_ (.A(_12663_),
    .X(_15014_));
 sky130_fd_sc_hd__and2_1 _19957_ (.A(_15014_),
    .B(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__and2_1 _19958_ (.A(_15014_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__and2_1 _19959_ (.A(_15014_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__and2_1 _19960_ (.A(_15014_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__and2_1 _19961_ (.A(_15014_),
    .B(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__and2_1 _19962_ (.A(_15014_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__buf_1 _19963_ (.A(_12663_),
    .X(_15015_));
 sky130_fd_sc_hd__and2_1 _19964_ (.A(_15015_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__and2_1 _19965_ (.A(_15015_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__and2_1 _19966_ (.A(_15015_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__and2_1 _19967_ (.A(_15015_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__and2_1 _19968_ (.A(_15015_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and2_1 _19969_ (.A(_15015_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_1 _19970_ (.A(_14536_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__and2_1 _19971_ (.A(_14536_),
    .B(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__xor2_1 _19972_ (.A(_02590_),
    .B(\decoded_imm_uj[1] ),
    .X(_01557_));
 sky130_fd_sc_hd__and2_1 _19973_ (.A(_02590_),
    .B(\decoded_imm_uj[1] ),
    .X(_15016_));
 sky130_fd_sc_hd__xnor2_1 _19974_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .Y(_15017_));
 sky130_fd_sc_hd__xnor2_1 _19975_ (.A(_15016_),
    .B(_15017_),
    .Y(_01562_));
 sky130_fd_sc_hd__xor2_1 _19976_ (.A(_01561_),
    .B(_02410_),
    .X(_01565_));
 sky130_fd_sc_hd__xor2_1 _19977_ (.A(_13247_),
    .B(_13250_),
    .X(_01567_));
 sky130_fd_sc_hd__xor2_1 _19978_ (.A(_13247_),
    .B(\decoded_imm_uj[3] ),
    .X(_15018_));
 sky130_fd_sc_hd__nand3b_2 _19979_ (.A_N(_15017_),
    .B(_02590_),
    .C(\decoded_imm_uj[1] ),
    .Y(_15019_));
 sky130_fd_sc_hd__nand2_1 _19980_ (.A(_13250_),
    .B(\decoded_imm_uj[2] ),
    .Y(_15020_));
 sky130_fd_sc_hd__nand2_1 _19981_ (.A(_15019_),
    .B(_15020_),
    .Y(_15021_));
 sky130_fd_sc_hd__xor2_1 _19982_ (.A(_15018_),
    .B(_15021_),
    .X(_01568_));
 sky130_fd_sc_hd__and2_1 _19983_ (.A(_13247_),
    .B(_13250_),
    .X(_15022_));
 sky130_fd_sc_hd__xor2_1 _19984_ (.A(_02582_),
    .B(_15022_),
    .X(_01571_));
 sky130_fd_sc_hd__xnor2_1 _19985_ (.A(\decoded_imm_uj[4] ),
    .B(_01475_),
    .Y(_15023_));
 sky130_fd_sc_hd__a2bb2oi_1 _19986_ (.A1_N(_02571_),
    .A2_N(\decoded_imm_uj[3] ),
    .B1(_15020_),
    .B2(_15019_),
    .Y(_15024_));
 sky130_fd_sc_hd__a21o_1 _19987_ (.A1(_02571_),
    .A2(\decoded_imm_uj[3] ),
    .B1(_15024_),
    .X(_15025_));
 sky130_fd_sc_hd__xor2_1 _19988_ (.A(_15023_),
    .B(_15025_),
    .X(_01572_));
 sky130_fd_sc_hd__clkbuf_2 _19989_ (.A(_02583_),
    .X(_15026_));
 sky130_fd_sc_hd__and3b_1 _19990_ (.A_N(_01475_),
    .B(_13247_),
    .C(_13250_),
    .X(_15027_));
 sky130_fd_sc_hd__xor2_1 _19991_ (.A(_15026_),
    .B(_15027_),
    .X(_01575_));
 sky130_fd_sc_hd__xor2_1 _19992_ (.A(_15026_),
    .B(\decoded_imm_uj[5] ),
    .X(_15028_));
 sky130_fd_sc_hd__o21ai_1 _19993_ (.A1(\decoded_imm_uj[4] ),
    .A2(_02582_),
    .B1(_15025_),
    .Y(_15029_));
 sky130_fd_sc_hd__o21ai_1 _19994_ (.A1(_00367_),
    .A2(_01475_),
    .B1(_15029_),
    .Y(_15030_));
 sky130_fd_sc_hd__xor2_1 _19995_ (.A(_15028_),
    .B(_15030_),
    .X(_01576_));
 sky130_fd_sc_hd__and4_1 _19996_ (.A(_02582_),
    .B(_15026_),
    .C(_13247_),
    .D(_13250_),
    .X(_15031_));
 sky130_fd_sc_hd__xor2_1 _19997_ (.A(_13239_),
    .B(_15031_),
    .X(_01579_));
 sky130_fd_sc_hd__nor2_1 _19998_ (.A(_13239_),
    .B(\decoded_imm_uj[6] ),
    .Y(_15032_));
 sky130_fd_sc_hd__and2_1 _19999_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .X(_15033_));
 sky130_fd_sc_hd__nor2_1 _20000_ (.A(_15032_),
    .B(_15033_),
    .Y(_15034_));
 sky130_fd_sc_hd__o21ai_1 _20001_ (.A1(_15026_),
    .A2(\decoded_imm_uj[5] ),
    .B1(_15030_),
    .Y(_15035_));
 sky130_fd_sc_hd__o21ai_2 _20002_ (.A1(_13242_),
    .A2(_14560_),
    .B1(_15035_),
    .Y(_15036_));
 sky130_fd_sc_hd__xor2_1 _20003_ (.A(_15034_),
    .B(_15036_),
    .X(_01580_));
 sky130_fd_sc_hd__clkbuf_2 _20004_ (.A(_02585_),
    .X(_15037_));
 sky130_fd_sc_hd__and4_1 _20005_ (.A(_15022_),
    .B(_13239_),
    .C(_15026_),
    .D(_02582_),
    .X(_15038_));
 sky130_fd_sc_hd__xor2_1 _20006_ (.A(_15037_),
    .B(_15038_),
    .X(_01583_));
 sky130_fd_sc_hd__xor2_1 _20007_ (.A(_15037_),
    .B(\decoded_imm_uj[7] ),
    .X(_15039_));
 sky130_vsdinv _20008_ (.A(_15032_),
    .Y(_15040_));
 sky130_fd_sc_hd__a21o_1 _20009_ (.A1(_15036_),
    .A2(_15040_),
    .B1(_15033_),
    .X(_15041_));
 sky130_fd_sc_hd__xor2_1 _20010_ (.A(_15039_),
    .B(_15041_),
    .X(_01584_));
 sky130_fd_sc_hd__and4_1 _20011_ (.A(_15027_),
    .B(_15037_),
    .C(_13239_),
    .D(_15026_),
    .X(_15042_));
 sky130_fd_sc_hd__xor2_1 _20012_ (.A(_13232_),
    .B(_15042_),
    .X(_01587_));
 sky130_fd_sc_hd__nor2_1 _20013_ (.A(_13232_),
    .B(\decoded_imm_uj[8] ),
    .Y(_15043_));
 sky130_fd_sc_hd__and2_1 _20014_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .X(_15044_));
 sky130_fd_sc_hd__nor2_1 _20015_ (.A(_15043_),
    .B(_15044_),
    .Y(_15045_));
 sky130_fd_sc_hd__o21ai_1 _20016_ (.A1(_15037_),
    .A2(\decoded_imm_uj[7] ),
    .B1(_15041_),
    .Y(_15046_));
 sky130_fd_sc_hd__o21ai_2 _20017_ (.A1(_13235_),
    .A2(_14564_),
    .B1(_15046_),
    .Y(_15047_));
 sky130_fd_sc_hd__xor2_1 _20018_ (.A(_15045_),
    .B(_15047_),
    .X(_01588_));
 sky130_fd_sc_hd__and4_1 _20019_ (.A(_15031_),
    .B(_13232_),
    .C(_15037_),
    .D(_13239_),
    .X(_15048_));
 sky130_fd_sc_hd__xor2_1 _20020_ (.A(_13230_),
    .B(_15048_),
    .X(_01591_));
 sky130_fd_sc_hd__xor2_1 _20021_ (.A(_13230_),
    .B(\decoded_imm_uj[9] ),
    .X(_15049_));
 sky130_vsdinv _20022_ (.A(_15043_),
    .Y(_15050_));
 sky130_fd_sc_hd__a21o_1 _20023_ (.A1(_15047_),
    .A2(_15050_),
    .B1(_15044_),
    .X(_15051_));
 sky130_fd_sc_hd__xor2_1 _20024_ (.A(_15049_),
    .B(_15051_),
    .X(_01592_));
 sky130_fd_sc_hd__and4_1 _20025_ (.A(_15038_),
    .B(_13230_),
    .C(_13232_),
    .D(_15037_),
    .X(_15052_));
 sky130_fd_sc_hd__xor2_1 _20026_ (.A(_13227_),
    .B(_15052_),
    .X(_01595_));
 sky130_fd_sc_hd__nor2_1 _20027_ (.A(_13227_),
    .B(\decoded_imm_uj[10] ),
    .Y(_15053_));
 sky130_fd_sc_hd__and2_1 _20028_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .X(_15054_));
 sky130_fd_sc_hd__nor2_1 _20029_ (.A(_15053_),
    .B(_15054_),
    .Y(_15055_));
 sky130_fd_sc_hd__or2_1 _20030_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .X(_15056_));
 sky130_fd_sc_hd__and2_1 _20031_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .X(_15057_));
 sky130_fd_sc_hd__a21o_1 _20032_ (.A1(_15051_),
    .A2(_15056_),
    .B1(_15057_),
    .X(_15058_));
 sky130_fd_sc_hd__xor2_1 _20033_ (.A(_15055_),
    .B(_15058_),
    .X(_01596_));
 sky130_fd_sc_hd__and4_1 _20034_ (.A(_15042_),
    .B(_13227_),
    .C(_13230_),
    .D(_13232_),
    .X(_15059_));
 sky130_fd_sc_hd__xor2_1 _20035_ (.A(_13224_),
    .B(_15059_),
    .X(_01599_));
 sky130_fd_sc_hd__xor2_2 _20036_ (.A(_02589_),
    .B(\decoded_imm_uj[11] ),
    .X(_15060_));
 sky130_vsdinv _20037_ (.A(_15053_),
    .Y(_15061_));
 sky130_fd_sc_hd__a21o_1 _20038_ (.A1(_15058_),
    .A2(_15061_),
    .B1(_15054_),
    .X(_15062_));
 sky130_fd_sc_hd__xor2_1 _20039_ (.A(_15060_),
    .B(_15062_),
    .X(_01600_));
 sky130_fd_sc_hd__and4_1 _20040_ (.A(_15048_),
    .B(_13224_),
    .C(_13227_),
    .D(_13230_),
    .X(_15063_));
 sky130_fd_sc_hd__xor2_1 _20041_ (.A(_13218_),
    .B(_15063_),
    .X(_01603_));
 sky130_fd_sc_hd__nand2_1 _20042_ (.A(_15062_),
    .B(_15060_),
    .Y(_15064_));
 sky130_fd_sc_hd__nand2_1 _20043_ (.A(_13224_),
    .B(\decoded_imm_uj[11] ),
    .Y(_15065_));
 sky130_fd_sc_hd__xor2_1 _20044_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .X(_15066_));
 sky130_fd_sc_hd__a21boi_1 _20045_ (.A1(_15064_),
    .A2(_15065_),
    .B1_N(_15066_),
    .Y(_15067_));
 sky130_fd_sc_hd__and3b_1 _20046_ (.A_N(_15066_),
    .B(_15064_),
    .C(_15065_),
    .X(_15068_));
 sky130_fd_sc_hd__nor2_1 _20047_ (.A(_15067_),
    .B(_15068_),
    .Y(_01604_));
 sky130_fd_sc_hd__and4_1 _20048_ (.A(_15052_),
    .B(_13218_),
    .C(_13224_),
    .D(_13227_),
    .X(_15069_));
 sky130_fd_sc_hd__xor2_1 _20049_ (.A(_13216_),
    .B(_15069_),
    .X(_01607_));
 sky130_fd_sc_hd__xor2_2 _20050_ (.A(_02562_),
    .B(\decoded_imm_uj[13] ),
    .X(_15070_));
 sky130_fd_sc_hd__a21o_1 _20051_ (.A1(_13218_),
    .A2(\decoded_imm_uj[12] ),
    .B1(_15067_),
    .X(_15071_));
 sky130_fd_sc_hd__xor2_1 _20052_ (.A(_15070_),
    .B(_15071_),
    .X(_01608_));
 sky130_fd_sc_hd__and4_1 _20053_ (.A(_15059_),
    .B(_13216_),
    .C(_13218_),
    .D(_13224_),
    .X(_15072_));
 sky130_fd_sc_hd__xor2_1 _20054_ (.A(_02563_),
    .B(_15072_),
    .X(_01611_));
 sky130_fd_sc_hd__xor2_2 _20055_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .X(_15073_));
 sky130_fd_sc_hd__and2_1 _20056_ (.A(_13216_),
    .B(\decoded_imm_uj[13] ),
    .X(_15074_));
 sky130_fd_sc_hd__a21o_1 _20057_ (.A1(_15071_),
    .A2(_15070_),
    .B1(_15074_),
    .X(_15075_));
 sky130_fd_sc_hd__xor2_1 _20058_ (.A(_15073_),
    .B(_15075_),
    .X(_01612_));
 sky130_fd_sc_hd__and4_1 _20059_ (.A(_15063_),
    .B(_02563_),
    .C(_13216_),
    .D(_13218_),
    .X(_15076_));
 sky130_fd_sc_hd__xor2_1 _20060_ (.A(_13209_),
    .B(_15076_),
    .X(_01615_));
 sky130_fd_sc_hd__xor2_2 _20061_ (.A(_02564_),
    .B(\decoded_imm_uj[15] ),
    .X(_15077_));
 sky130_fd_sc_hd__nand2_1 _20062_ (.A(_15075_),
    .B(_15073_),
    .Y(_15078_));
 sky130_fd_sc_hd__o21ai_2 _20063_ (.A1(_13212_),
    .A2(_14586_),
    .B1(_15078_),
    .Y(_15079_));
 sky130_fd_sc_hd__xor2_1 _20064_ (.A(_15077_),
    .B(_15079_),
    .X(_01616_));
 sky130_fd_sc_hd__and4_1 _20065_ (.A(_15069_),
    .B(_13209_),
    .C(_02563_),
    .D(_13216_),
    .X(_15080_));
 sky130_fd_sc_hd__xor2_1 _20066_ (.A(_13206_),
    .B(_15080_),
    .X(_01619_));
 sky130_fd_sc_hd__xor2_2 _20067_ (.A(_02565_),
    .B(\decoded_imm_uj[16] ),
    .X(_15081_));
 sky130_fd_sc_hd__and2_1 _20068_ (.A(_15079_),
    .B(_15077_),
    .X(_15082_));
 sky130_fd_sc_hd__a21o_1 _20069_ (.A1(_13209_),
    .A2(\decoded_imm_uj[15] ),
    .B1(_15082_),
    .X(_15083_));
 sky130_fd_sc_hd__xor2_1 _20070_ (.A(_15081_),
    .B(_15083_),
    .X(_01620_));
 sky130_fd_sc_hd__and4_1 _20071_ (.A(_15072_),
    .B(_13206_),
    .C(_13209_),
    .D(_02563_),
    .X(_15084_));
 sky130_fd_sc_hd__xor2_1 _20072_ (.A(_13202_),
    .B(_15084_),
    .X(_01623_));
 sky130_fd_sc_hd__xor2_2 _20073_ (.A(_02566_),
    .B(\decoded_imm_uj[17] ),
    .X(_15085_));
 sky130_fd_sc_hd__and2_1 _20074_ (.A(_13206_),
    .B(\decoded_imm_uj[16] ),
    .X(_15086_));
 sky130_fd_sc_hd__a21o_1 _20075_ (.A1(_15083_),
    .A2(_15081_),
    .B1(_15086_),
    .X(_15087_));
 sky130_fd_sc_hd__xor2_1 _20076_ (.A(_15085_),
    .B(_15087_),
    .X(_01624_));
 sky130_fd_sc_hd__and4_1 _20077_ (.A(_15076_),
    .B(_13202_),
    .C(_13206_),
    .D(_13209_),
    .X(_15088_));
 sky130_fd_sc_hd__xor2_1 _20078_ (.A(_13200_),
    .B(_15088_),
    .X(_01627_));
 sky130_fd_sc_hd__nor2_1 _20079_ (.A(_13200_),
    .B(\decoded_imm_uj[18] ),
    .Y(_15089_));
 sky130_fd_sc_hd__and2_1 _20080_ (.A(_02567_),
    .B(\decoded_imm_uj[18] ),
    .X(_15090_));
 sky130_fd_sc_hd__nor2_1 _20081_ (.A(_15089_),
    .B(_15090_),
    .Y(_15091_));
 sky130_fd_sc_hd__and2_1 _20082_ (.A(_13202_),
    .B(\decoded_imm_uj[17] ),
    .X(_15092_));
 sky130_fd_sc_hd__a21o_1 _20083_ (.A1(_15087_),
    .A2(_15085_),
    .B1(_15092_),
    .X(_15093_));
 sky130_fd_sc_hd__xor2_1 _20084_ (.A(_15091_),
    .B(_15093_),
    .X(_01628_));
 sky130_fd_sc_hd__and4_1 _20085_ (.A(_15080_),
    .B(_13200_),
    .C(_13202_),
    .D(_13206_),
    .X(_15094_));
 sky130_fd_sc_hd__xor2_1 _20086_ (.A(_13197_),
    .B(_15094_),
    .X(_01631_));
 sky130_fd_sc_hd__xor2_4 _20087_ (.A(_02568_),
    .B(\decoded_imm_uj[19] ),
    .X(_15095_));
 sky130_vsdinv _20088_ (.A(_15089_),
    .Y(_15096_));
 sky130_fd_sc_hd__a21o_1 _20089_ (.A1(_15093_),
    .A2(_15096_),
    .B1(_15090_),
    .X(_15097_));
 sky130_fd_sc_hd__xor2_1 _20090_ (.A(_15095_),
    .B(_15097_),
    .X(_01632_));
 sky130_fd_sc_hd__and4_1 _20091_ (.A(_15084_),
    .B(_13197_),
    .C(_13200_),
    .D(_13202_),
    .X(_15098_));
 sky130_fd_sc_hd__xor2_1 _20092_ (.A(_02569_),
    .B(_15098_),
    .X(_01635_));
 sky130_fd_sc_hd__xnor2_1 _20093_ (.A(_02569_),
    .B(_14127_),
    .Y(_15099_));
 sky130_fd_sc_hd__and2_1 _20094_ (.A(_13197_),
    .B(\decoded_imm_uj[19] ),
    .X(_15100_));
 sky130_fd_sc_hd__a21oi_2 _20095_ (.A1(_15097_),
    .A2(_15095_),
    .B1(_15100_),
    .Y(_15101_));
 sky130_fd_sc_hd__xor2_1 _20096_ (.A(_15099_),
    .B(_15101_),
    .X(_01636_));
 sky130_fd_sc_hd__and4_1 _20097_ (.A(_15088_),
    .B(_02569_),
    .C(_13197_),
    .D(_13200_),
    .X(_15102_));
 sky130_fd_sc_hd__xor2_1 _20098_ (.A(_13188_),
    .B(_15102_),
    .X(_01639_));
 sky130_fd_sc_hd__xor2_4 _20099_ (.A(_02570_),
    .B(\decoded_imm_uj[20] ),
    .X(_15103_));
 sky130_fd_sc_hd__a21o_1 _20100_ (.A1(_13191_),
    .A2(_14630_),
    .B1(_15101_),
    .X(_15104_));
 sky130_fd_sc_hd__o21ai_2 _20101_ (.A1(_13191_),
    .A2(_14630_),
    .B1(_15104_),
    .Y(_15105_));
 sky130_fd_sc_hd__xor2_1 _20102_ (.A(_15103_),
    .B(_15105_),
    .X(_01640_));
 sky130_fd_sc_hd__and4_1 _20103_ (.A(_15094_),
    .B(_13188_),
    .C(_02569_),
    .D(_13197_),
    .X(_15106_));
 sky130_fd_sc_hd__xor2_1 _20104_ (.A(_13185_),
    .B(_15106_),
    .X(_01643_));
 sky130_fd_sc_hd__xor2_4 _20105_ (.A(_02572_),
    .B(_14124_),
    .X(_15107_));
 sky130_fd_sc_hd__and2_1 _20106_ (.A(_13188_),
    .B(_14125_),
    .X(_15108_));
 sky130_fd_sc_hd__a21oi_1 _20107_ (.A1(_15105_),
    .A2(_15103_),
    .B1(_15108_),
    .Y(_15109_));
 sky130_fd_sc_hd__xnor2_1 _20108_ (.A(_15107_),
    .B(_15109_),
    .Y(_01644_));
 sky130_fd_sc_hd__and4_1 _20109_ (.A(_15098_),
    .B(_02572_),
    .C(_02570_),
    .D(_02569_),
    .X(_15110_));
 sky130_fd_sc_hd__xor2_1 _20110_ (.A(_13183_),
    .B(_15110_),
    .X(_01647_));
 sky130_fd_sc_hd__xor2_4 _20111_ (.A(_02573_),
    .B(_14124_),
    .X(_15111_));
 sky130_fd_sc_hd__and2_1 _20112_ (.A(_13185_),
    .B(_14126_),
    .X(_15112_));
 sky130_fd_sc_hd__a311o_1 _20113_ (.A1(_15105_),
    .A2(_15103_),
    .A3(_15107_),
    .B1(_15108_),
    .C1(_15112_),
    .X(_15113_));
 sky130_fd_sc_hd__xor2_1 _20114_ (.A(_15111_),
    .B(_15113_),
    .X(_01648_));
 sky130_fd_sc_hd__and4_1 _20115_ (.A(_15102_),
    .B(_13183_),
    .C(_13185_),
    .D(_13188_),
    .X(_15114_));
 sky130_fd_sc_hd__xor2_1 _20116_ (.A(_13179_),
    .B(_15114_),
    .X(_01651_));
 sky130_fd_sc_hd__xor2_2 _20117_ (.A(_02574_),
    .B(_14124_),
    .X(_15115_));
 sky130_fd_sc_hd__and2_1 _20118_ (.A(_13183_),
    .B(_14127_),
    .X(_15116_));
 sky130_fd_sc_hd__a21oi_1 _20119_ (.A1(_15113_),
    .A2(_15111_),
    .B1(_15116_),
    .Y(_15117_));
 sky130_fd_sc_hd__xnor2_1 _20120_ (.A(_15115_),
    .B(_15117_),
    .Y(_01652_));
 sky130_fd_sc_hd__and4_1 _20121_ (.A(_15106_),
    .B(_13179_),
    .C(_13183_),
    .D(_13185_),
    .X(_15118_));
 sky130_fd_sc_hd__xor2_1 _20122_ (.A(_13176_),
    .B(_15118_),
    .X(_01655_));
 sky130_fd_sc_hd__xor2_4 _20123_ (.A(_02575_),
    .B(_14124_),
    .X(_15119_));
 sky130_fd_sc_hd__nand3_1 _20124_ (.A(_15105_),
    .B(_15103_),
    .C(_15107_),
    .Y(_15120_));
 sky130_fd_sc_hd__nand3b_1 _20125_ (.A_N(_15120_),
    .B(_15111_),
    .C(_15115_),
    .Y(_15121_));
 sky130_fd_sc_hd__o41ai_2 _20126_ (.A1(_13179_),
    .A2(_02573_),
    .A3(_13185_),
    .A4(_13188_),
    .B1(_14124_),
    .Y(_15122_));
 sky130_fd_sc_hd__nand2_2 _20127_ (.A(_15121_),
    .B(_15122_),
    .Y(_15123_));
 sky130_fd_sc_hd__xor2_1 _20128_ (.A(_15119_),
    .B(_15123_),
    .X(_01656_));
 sky130_fd_sc_hd__and4_1 _20129_ (.A(_15110_),
    .B(_13176_),
    .C(_13179_),
    .D(_13183_),
    .X(_15124_));
 sky130_fd_sc_hd__xor2_1 _20130_ (.A(_02576_),
    .B(_15124_),
    .X(_01659_));
 sky130_fd_sc_hd__xor2_2 _20131_ (.A(_02576_),
    .B(_14125_),
    .X(_15125_));
 sky130_fd_sc_hd__and2_1 _20132_ (.A(_13176_),
    .B(_14125_),
    .X(_15126_));
 sky130_fd_sc_hd__a21oi_1 _20133_ (.A1(_15123_),
    .A2(_15119_),
    .B1(_15126_),
    .Y(_15127_));
 sky130_fd_sc_hd__xnor2_1 _20134_ (.A(_15125_),
    .B(_15127_),
    .Y(_01660_));
 sky130_fd_sc_hd__and4_1 _20135_ (.A(_15114_),
    .B(_02576_),
    .C(_13176_),
    .D(_13179_),
    .X(_15128_));
 sky130_fd_sc_hd__xor2_1 _20136_ (.A(_13167_),
    .B(_15128_),
    .X(_01663_));
 sky130_fd_sc_hd__xor2_4 _20137_ (.A(_02577_),
    .B(_14125_),
    .X(_15129_));
 sky130_vsdinv _20138_ (.A(_15126_),
    .Y(_15130_));
 sky130_fd_sc_hd__nand3_2 _20139_ (.A(_15123_),
    .B(_15119_),
    .C(_15125_),
    .Y(_15131_));
 sky130_fd_sc_hd__o211ai_2 _20140_ (.A1(_13172_),
    .A2(_14630_),
    .B1(_15130_),
    .C1(_15131_),
    .Y(_15132_));
 sky130_fd_sc_hd__xor2_1 _20141_ (.A(_15129_),
    .B(_15132_),
    .X(_01664_));
 sky130_fd_sc_hd__and4_1 _20142_ (.A(_15118_),
    .B(_13167_),
    .C(_02576_),
    .D(_13176_),
    .X(_15133_));
 sky130_fd_sc_hd__xor2_1 _20143_ (.A(_02578_),
    .B(_15133_),
    .X(_01667_));
 sky130_fd_sc_hd__xor2_2 _20144_ (.A(_02578_),
    .B(_14125_),
    .X(_15134_));
 sky130_fd_sc_hd__and2_1 _20145_ (.A(_13167_),
    .B(_14127_),
    .X(_15135_));
 sky130_fd_sc_hd__a21oi_1 _20146_ (.A1(_15132_),
    .A2(_15129_),
    .B1(_15135_),
    .Y(_15136_));
 sky130_fd_sc_hd__xnor2_1 _20147_ (.A(_15134_),
    .B(_15136_),
    .Y(_01668_));
 sky130_fd_sc_hd__and4_1 _20148_ (.A(_15124_),
    .B(_02578_),
    .C(_13167_),
    .D(_02576_),
    .X(_15137_));
 sky130_fd_sc_hd__xor2_1 _20149_ (.A(_13160_),
    .B(_15137_),
    .X(_01671_));
 sky130_fd_sc_hd__xor2_4 _20150_ (.A(_02579_),
    .B(_14126_),
    .X(_15138_));
 sky130_fd_sc_hd__nand2_1 _20151_ (.A(_15129_),
    .B(_15134_),
    .Y(_15139_));
 sky130_fd_sc_hd__a41oi_1 _20152_ (.A1(_13164_),
    .A2(_13168_),
    .A3(_13172_),
    .A4(_13177_),
    .B1(_14630_),
    .Y(_15140_));
 sky130_fd_sc_hd__o21bai_2 _20153_ (.A1(_15139_),
    .A2(_15131_),
    .B1_N(_15140_),
    .Y(_15141_));
 sky130_fd_sc_hd__xor2_1 _20154_ (.A(_15138_),
    .B(_15141_),
    .X(_01672_));
 sky130_fd_sc_hd__and4_1 _20155_ (.A(_15128_),
    .B(_13160_),
    .C(_02578_),
    .D(_13167_),
    .X(_15142_));
 sky130_fd_sc_hd__xor2_1 _20156_ (.A(_02580_),
    .B(_15142_),
    .X(_01675_));
 sky130_fd_sc_hd__nand2_1 _20157_ (.A(_15141_),
    .B(_15138_),
    .Y(_15143_));
 sky130_fd_sc_hd__and2_1 _20158_ (.A(_13160_),
    .B(_14126_),
    .X(_15144_));
 sky130_vsdinv _20159_ (.A(_15144_),
    .Y(_15145_));
 sky130_fd_sc_hd__xnor2_1 _20160_ (.A(_02580_),
    .B(_14127_),
    .Y(_15146_));
 sky130_fd_sc_hd__a21oi_1 _20161_ (.A1(_15143_),
    .A2(_15145_),
    .B1(_15146_),
    .Y(_15147_));
 sky130_fd_sc_hd__and3_1 _20162_ (.A(_15143_),
    .B(_15145_),
    .C(_15146_),
    .X(_15148_));
 sky130_fd_sc_hd__nor2_1 _20163_ (.A(_15147_),
    .B(_15148_),
    .Y(_01676_));
 sky130_fd_sc_hd__nand3_1 _20164_ (.A(_15137_),
    .B(_02580_),
    .C(_13160_),
    .Y(_15149_));
 sky130_fd_sc_hd__xnor2_1 _20165_ (.A(_02581_),
    .B(_15149_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_1 _20166_ (.A(_13157_),
    .B(_14630_),
    .Y(_15150_));
 sky130_fd_sc_hd__nand3_1 _20167_ (.A(_15141_),
    .B(_15138_),
    .C(_15150_),
    .Y(_15151_));
 sky130_fd_sc_hd__o21ai_1 _20168_ (.A1(_02580_),
    .A2(_13160_),
    .B1(_14127_),
    .Y(_15152_));
 sky130_fd_sc_hd__xnor2_1 _20169_ (.A(_02581_),
    .B(_14126_),
    .Y(_15153_));
 sky130_fd_sc_hd__a21oi_1 _20170_ (.A1(_15151_),
    .A2(_15152_),
    .B1(_15153_),
    .Y(_15154_));
 sky130_fd_sc_hd__and3_1 _20171_ (.A(_15151_),
    .B(_15152_),
    .C(_15153_),
    .X(_15155_));
 sky130_fd_sc_hd__nor2_1 _20172_ (.A(_15154_),
    .B(_15155_),
    .Y(_01680_));
 sky130_fd_sc_hd__nor2_4 _20173_ (.A(_14658_),
    .B(\mem_wordsize[1] ),
    .Y(_01683_));
 sky130_vsdinv _20174_ (.A(_14264_),
    .Y(_15156_));
 sky130_fd_sc_hd__clkbuf_4 _20175_ (.A(_14658_),
    .X(_15157_));
 sky130_fd_sc_hd__a21o_1 _20176_ (.A1(_15156_),
    .A2(_15157_),
    .B1(_01683_),
    .X(_15158_));
 sky130_fd_sc_hd__o21a_1 _20177_ (.A1(_00304_),
    .A2(_15158_),
    .B1(net232),
    .X(_01684_));
 sky130_fd_sc_hd__nand3_1 _20178_ (.A(_00301_),
    .B(_14715_),
    .C(_01685_),
    .Y(_15159_));
 sky130_vsdinv _20179_ (.A(_15159_),
    .Y(_01686_));
 sky130_fd_sc_hd__and2b_1 _20180_ (.A_N(_14828_),
    .B(_14268_),
    .X(_15160_));
 sky130_fd_sc_hd__o21a_1 _20181_ (.A1(_15160_),
    .A2(_15158_),
    .B1(net232),
    .X(_01687_));
 sky130_fd_sc_hd__nand3_1 _20182_ (.A(_00301_),
    .B(_14715_),
    .C(_01688_),
    .Y(_15161_));
 sky130_vsdinv _20183_ (.A(_15161_),
    .Y(_01689_));
 sky130_fd_sc_hd__and2b_1 _20184_ (.A_N(_14267_),
    .B(_14263_),
    .X(_15162_));
 sky130_fd_sc_hd__a211o_4 _20185_ (.A1(_14828_),
    .A2(_15157_),
    .B1(net453),
    .C1(_15162_),
    .X(net235));
 sky130_fd_sc_hd__and2_1 _20186_ (.A(net235),
    .B(net232),
    .X(_01690_));
 sky130_fd_sc_hd__nand3_1 _20187_ (.A(_00301_),
    .B(_14715_),
    .C(_01691_),
    .Y(_15163_));
 sky130_vsdinv _20188_ (.A(_15163_),
    .Y(_01692_));
 sky130_fd_sc_hd__clkbuf_2 _20189_ (.A(_14267_),
    .X(_15164_));
 sky130_fd_sc_hd__and2_1 _20190_ (.A(_14264_),
    .B(_14658_),
    .X(_15165_));
 sky130_fd_sc_hd__a211o_4 _20191_ (.A1(_14828_),
    .A2(_15164_),
    .B1(net453),
    .C1(_15165_),
    .X(net236));
 sky130_fd_sc_hd__and2_1 _20192_ (.A(net236),
    .B(net232),
    .X(_01693_));
 sky130_fd_sc_hd__nand3_1 _20193_ (.A(_12670_),
    .B(_14715_),
    .C(_01694_),
    .Y(_15166_));
 sky130_vsdinv _20194_ (.A(_15166_),
    .Y(_01695_));
 sky130_fd_sc_hd__nor2_4 _20195_ (.A(\irq_pending[1] ),
    .B(net12),
    .Y(_01696_));
 sky130_fd_sc_hd__inv_2 _20196_ (.A(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__o21a_1 _20197_ (.A1(\irq_pending[1] ),
    .A2(net12),
    .B1(_13540_),
    .X(_01698_));
 sky130_fd_sc_hd__buf_6 _20198_ (.A(_12885_),
    .X(_15167_));
 sky130_fd_sc_hd__nand3_2 _20199_ (.A(_00297_),
    .B(_14634_),
    .C(_12893_),
    .Y(_15168_));
 sky130_fd_sc_hd__nor2_1 _20200_ (.A(_15167_),
    .B(_15168_),
    .Y(_01700_));
 sky130_fd_sc_hd__o21a_1 _20201_ (.A1(_14651_),
    .A2(_13540_),
    .B1(_01696_),
    .X(_01701_));
 sky130_fd_sc_hd__o2bb2ai_1 _20202_ (.A1_N(_01697_),
    .A2_N(_15168_),
    .B1(_14638_),
    .B2(_01704_),
    .Y(_01705_));
 sky130_vsdinv _20203_ (.A(net33),
    .Y(_01707_));
 sky130_fd_sc_hd__clkbuf_2 _20204_ (.A(_14828_),
    .X(_15169_));
 sky130_vsdinv _20205_ (.A(net306),
    .Y(_15170_));
 sky130_fd_sc_hd__clkbuf_2 _20206_ (.A(_15170_),
    .X(_15171_));
 sky130_vsdinv _20207_ (.A(net63),
    .Y(_01812_));
 sky130_fd_sc_hd__buf_4 _20208_ (.A(_14264_),
    .X(_15172_));
 sky130_fd_sc_hd__nand3b_1 _20209_ (.A_N(_15164_),
    .B(_15172_),
    .C(net40),
    .Y(_15173_));
 sky130_fd_sc_hd__nand3_1 _20210_ (.A(_14265_),
    .B(_14269_),
    .C(net49),
    .Y(_15174_));
 sky130_fd_sc_hd__o311a_1 _20211_ (.A1(_15169_),
    .A2(_15171_),
    .A3(_01812_),
    .B1(_15173_),
    .C1(_15174_),
    .X(_01708_));
 sky130_fd_sc_hd__clkbuf_4 _20212_ (.A(_15157_),
    .X(_15175_));
 sky130_fd_sc_hd__clkbuf_2 _20213_ (.A(_15175_),
    .X(_15176_));
 sky130_fd_sc_hd__clkbuf_2 _20214_ (.A(_14833_),
    .X(_15177_));
 sky130_fd_sc_hd__o2bb2a_1 _20215_ (.A1_N(_15176_),
    .A2_N(_01710_),
    .B1(_01709_),
    .B2(_15177_),
    .X(_01711_));
 sky130_fd_sc_hd__clkbuf_4 _20216_ (.A(_14182_),
    .X(_15178_));
 sky130_fd_sc_hd__and2_1 _20217_ (.A(\count_instr[32] ),
    .B(_14170_),
    .X(_15179_));
 sky130_fd_sc_hd__a221oi_2 _20218_ (.A1(\count_instr[0] ),
    .A2(_15178_),
    .B1(_14186_),
    .B2(\count_cycle[32] ),
    .C1(_15179_),
    .Y(_01715_));
 sky130_fd_sc_hd__nor3b_4 _20219_ (.A(_12830_),
    .B(_12907_),
    .C_N(_00370_),
    .Y(_15180_));
 sky130_fd_sc_hd__a221oi_2 _20220_ (.A1(\irq_mask[0] ),
    .A2(_14155_),
    .B1(_14138_),
    .B2(\timer[0] ),
    .C1(_15180_),
    .Y(_01718_));
 sky130_fd_sc_hd__buf_4 _20221_ (.A(_12659_),
    .X(_15181_));
 sky130_fd_sc_hd__clkbuf_4 _20222_ (.A(_12812_),
    .X(_15182_));
 sky130_fd_sc_hd__xnor2_1 _20223_ (.A(\decoded_imm[0] ),
    .B(\reg_next_pc[0] ),
    .Y(_15183_));
 sky130_fd_sc_hd__buf_4 _20224_ (.A(_13872_),
    .X(_15184_));
 sky130_fd_sc_hd__a2bb2oi_2 _20225_ (.A1_N(_01719_),
    .A2_N(_15184_),
    .B1(_14827_),
    .B2(_01713_),
    .Y(_15185_));
 sky130_fd_sc_hd__o221ai_2 _20226_ (.A1(_15181_),
    .A2(_01712_),
    .B1(_15182_),
    .B2(_15183_),
    .C1(_15185_),
    .Y(_01720_));
 sky130_vsdinv _20227_ (.A(net44),
    .Y(_01721_));
 sky130_vsdinv _20228_ (.A(net64),
    .Y(_01826_));
 sky130_fd_sc_hd__clkbuf_2 _20229_ (.A(_14264_),
    .X(_15186_));
 sky130_fd_sc_hd__nand3b_1 _20230_ (.A_N(_15164_),
    .B(_15186_),
    .C(net499),
    .Y(_15187_));
 sky130_fd_sc_hd__nand3_1 _20231_ (.A(_14265_),
    .B(_14269_),
    .C(net50),
    .Y(_15188_));
 sky130_fd_sc_hd__o311a_1 _20232_ (.A1(_15169_),
    .A2(_15171_),
    .A3(_01826_),
    .B1(_15187_),
    .C1(_15188_),
    .X(_01722_));
 sky130_fd_sc_hd__o2bb2a_1 _20233_ (.A1_N(_15176_),
    .A2_N(_01724_),
    .B1(_01723_),
    .B2(_15177_),
    .X(_01725_));
 sky130_vsdinv _20234_ (.A(\count_cycle[1] ),
    .Y(_01728_));
 sky130_fd_sc_hd__and2_1 _20235_ (.A(\count_instr[33] ),
    .B(_14170_),
    .X(_15189_));
 sky130_fd_sc_hd__a221oi_2 _20236_ (.A1(\count_instr[1] ),
    .A2(_15178_),
    .B1(_14186_),
    .B2(\count_cycle[33] ),
    .C1(_15189_),
    .Y(_01729_));
 sky130_fd_sc_hd__nand2_4 _20237_ (.A(_12830_),
    .B(_12831_),
    .Y(_15190_));
 sky130_fd_sc_hd__clkbuf_4 _20238_ (.A(_15190_),
    .X(_15191_));
 sky130_fd_sc_hd__and2_1 _20239_ (.A(_13540_),
    .B(_12955_),
    .X(_15192_));
 sky130_fd_sc_hd__a221oi_2 _20240_ (.A1(_14139_),
    .A2(\timer[1] ),
    .B1(\cpuregs_rs1[1] ),
    .B2(_15191_),
    .C1(_15192_),
    .Y(_01731_));
 sky130_fd_sc_hd__and2_1 _20241_ (.A(\decoded_imm[0] ),
    .B(\reg_next_pc[0] ),
    .X(_15193_));
 sky130_fd_sc_hd__xor2_4 _20242_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .X(_15194_));
 sky130_fd_sc_hd__xor2_2 _20243_ (.A(_15193_),
    .B(_15194_),
    .X(_15195_));
 sky130_fd_sc_hd__and2b_1 _20244_ (.A_N(_01726_),
    .B(_12652_),
    .X(_15196_));
 sky130_fd_sc_hd__buf_4 _20245_ (.A(_12853_),
    .X(_15197_));
 sky130_fd_sc_hd__o2bb2ai_2 _20246_ (.A1_N(_15167_),
    .A2_N(_01727_),
    .B1(_01732_),
    .B2(_15197_),
    .Y(_15198_));
 sky130_fd_sc_hd__a211o_1 _20247_ (.A1(_15195_),
    .A2(_14822_),
    .B1(_15196_),
    .C1(_15198_),
    .X(_01733_));
 sky130_vsdinv _20248_ (.A(net55),
    .Y(_01734_));
 sky130_vsdinv _20249_ (.A(net34),
    .Y(_01839_));
 sky130_fd_sc_hd__nand3b_1 _20250_ (.A_N(_15164_),
    .B(_15186_),
    .C(net42),
    .Y(_15199_));
 sky130_fd_sc_hd__nand3_1 _20251_ (.A(_14265_),
    .B(_14269_),
    .C(net51),
    .Y(_15200_));
 sky130_fd_sc_hd__o311a_1 _20252_ (.A1(_15169_),
    .A2(_15171_),
    .A3(_01839_),
    .B1(_15199_),
    .C1(_15200_),
    .X(_01735_));
 sky130_fd_sc_hd__clkbuf_2 _20253_ (.A(_14833_),
    .X(_15201_));
 sky130_fd_sc_hd__o2bb2a_1 _20254_ (.A1_N(_15176_),
    .A2_N(_01737_),
    .B1(_01736_),
    .B2(_15201_),
    .X(_01738_));
 sky130_fd_sc_hd__and2_1 _20255_ (.A(_14185_),
    .B(_13596_),
    .X(_15202_));
 sky130_fd_sc_hd__a221oi_2 _20256_ (.A1(\count_instr[34] ),
    .A2(_14171_),
    .B1(\count_instr[2] ),
    .B2(_14183_),
    .C1(_15202_),
    .Y(_01742_));
 sky130_fd_sc_hd__buf_1 _20257_ (.A(_12908_),
    .X(_15203_));
 sky130_fd_sc_hd__and2_1 _20258_ (.A(\irq_mask[2] ),
    .B(_15203_),
    .X(_15204_));
 sky130_fd_sc_hd__a221oi_2 _20259_ (.A1(_14139_),
    .A2(\timer[2] ),
    .B1(\cpuregs_rs1[2] ),
    .B2(_15191_),
    .C1(_15204_),
    .Y(_01744_));
 sky130_fd_sc_hd__buf_4 _20260_ (.A(_12659_),
    .X(_04073_));
 sky130_fd_sc_hd__nor2_1 _20261_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .Y(_04074_));
 sky130_fd_sc_hd__and2_1 _20262_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .X(_04075_));
 sky130_fd_sc_hd__nor2_2 _20263_ (.A(_04074_),
    .B(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__and2_1 _20264_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .X(_04077_));
 sky130_fd_sc_hd__a21o_1 _20265_ (.A1(_15194_),
    .A2(_15193_),
    .B1(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__xnor2_2 _20266_ (.A(_04076_),
    .B(_04078_),
    .Y(_04079_));
 sky130_fd_sc_hd__buf_6 _20267_ (.A(_12843_),
    .X(_04080_));
 sky130_fd_sc_hd__a2bb2oi_4 _20268_ (.A1_N(_01745_),
    .A2_N(_15184_),
    .B1(_04080_),
    .B2(_01740_),
    .Y(_04081_));
 sky130_fd_sc_hd__o221ai_4 _20269_ (.A1(_04073_),
    .A2(_01739_),
    .B1(_15182_),
    .B2(_04079_),
    .C1(_04081_),
    .Y(_01746_));
 sky130_vsdinv _20270_ (.A(net58),
    .Y(_01747_));
 sky130_vsdinv _20271_ (.A(net35),
    .Y(_01852_));
 sky130_fd_sc_hd__nand3b_1 _20272_ (.A_N(_15164_),
    .B(_15186_),
    .C(net498),
    .Y(_04082_));
 sky130_fd_sc_hd__nand3_1 _20273_ (.A(_15172_),
    .B(_14829_),
    .C(net52),
    .Y(_04083_));
 sky130_fd_sc_hd__o311a_1 _20274_ (.A1(_15169_),
    .A2(_15171_),
    .A3(_01852_),
    .B1(_04082_),
    .C1(_04083_),
    .X(_01748_));
 sky130_fd_sc_hd__o2bb2a_1 _20275_ (.A1_N(_15176_),
    .A2_N(_01750_),
    .B1(_01749_),
    .B2(_15201_),
    .X(_01751_));
 sky130_fd_sc_hd__and2_1 _20276_ (.A(\count_instr[35] ),
    .B(_14170_),
    .X(_04084_));
 sky130_fd_sc_hd__a221oi_2 _20277_ (.A1(\count_instr[3] ),
    .A2(_15178_),
    .B1(_14186_),
    .B2(\count_cycle[35] ),
    .C1(_04084_),
    .Y(_01755_));
 sky130_fd_sc_hd__buf_1 _20278_ (.A(net494),
    .X(_04085_));
 sky130_fd_sc_hd__and2_1 _20279_ (.A(_04085_),
    .B(\timer[3] ),
    .X(_04086_));
 sky130_fd_sc_hd__a221oi_2 _20280_ (.A1(\irq_mask[3] ),
    .A2(_14155_),
    .B1(\cpuregs_rs1[3] ),
    .B2(_15191_),
    .C1(_04086_),
    .Y(_01757_));
 sky130_fd_sc_hd__and2_1 _20281_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .X(_04087_));
 sky130_fd_sc_hd__nor2_2 _20282_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_04088_));
 sky130_vsdinv _20283_ (.A(_04074_),
    .Y(_04089_));
 sky130_fd_sc_hd__a21oi_4 _20284_ (.A1(_04078_),
    .A2(_04089_),
    .B1(_04075_),
    .Y(_04090_));
 sky130_fd_sc_hd__o21a_1 _20285_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__buf_4 _20286_ (.A(_12845_),
    .X(_04092_));
 sky130_fd_sc_hd__o31ai_1 _20287_ (.A1(_04087_),
    .A2(_04088_),
    .A3(_04090_),
    .B1(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__buf_6 _20288_ (.A(_13872_),
    .X(_04094_));
 sky130_fd_sc_hd__a2bb2oi_2 _20289_ (.A1_N(_01758_),
    .A2_N(_04094_),
    .B1(_04080_),
    .B2(_01753_),
    .Y(_04095_));
 sky130_fd_sc_hd__o221ai_1 _20290_ (.A1(_04073_),
    .A2(_01752_),
    .B1(_04091_),
    .B2(_04093_),
    .C1(_04095_),
    .Y(_01759_));
 sky130_vsdinv _20291_ (.A(net59),
    .Y(_01760_));
 sky130_vsdinv _20292_ (.A(net36),
    .Y(_01865_));
 sky130_fd_sc_hd__nand3b_1 _20293_ (.A_N(_15164_),
    .B(_15186_),
    .C(net45),
    .Y(_04096_));
 sky130_fd_sc_hd__nand3_1 _20294_ (.A(_15172_),
    .B(_14829_),
    .C(net53),
    .Y(_04097_));
 sky130_fd_sc_hd__o311a_1 _20295_ (.A1(_15169_),
    .A2(_15171_),
    .A3(_01865_),
    .B1(_04096_),
    .C1(_04097_),
    .X(_01761_));
 sky130_fd_sc_hd__clkbuf_4 _20296_ (.A(_15157_),
    .X(_04098_));
 sky130_fd_sc_hd__o2bb2a_1 _20297_ (.A1_N(_04098_),
    .A2_N(_01763_),
    .B1(_01762_),
    .B2(_15201_),
    .X(_01764_));
 sky130_fd_sc_hd__clkbuf_4 _20298_ (.A(_14182_),
    .X(_04099_));
 sky130_fd_sc_hd__and2_1 _20299_ (.A(\count_instr[36] ),
    .B(_14170_),
    .X(_04100_));
 sky130_fd_sc_hd__a221oi_2 _20300_ (.A1(\count_instr[4] ),
    .A2(_04099_),
    .B1(_14186_),
    .B2(\count_cycle[36] ),
    .C1(_04100_),
    .Y(_01768_));
 sky130_fd_sc_hd__and2_1 _20301_ (.A(_04085_),
    .B(\timer[4] ),
    .X(_04101_));
 sky130_fd_sc_hd__a221oi_2 _20302_ (.A1(\irq_mask[4] ),
    .A2(_14155_),
    .B1(\cpuregs_rs1[4] ),
    .B2(_15191_),
    .C1(_04101_),
    .Y(_01770_));
 sky130_fd_sc_hd__xor2_4 _20303_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .X(_04102_));
 sky130_fd_sc_hd__o21bai_2 _20304_ (.A1(_04088_),
    .A2(_04090_),
    .B1_N(_04087_),
    .Y(_04103_));
 sky130_fd_sc_hd__xnor2_1 _20305_ (.A(_04102_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__a2bb2oi_4 _20306_ (.A1_N(_01771_),
    .A2_N(_04094_),
    .B1(_04080_),
    .B2(_01766_),
    .Y(_04105_));
 sky130_fd_sc_hd__o221ai_2 _20307_ (.A1(_04073_),
    .A2(_01765_),
    .B1(_15182_),
    .B2(_04104_),
    .C1(_04105_),
    .Y(_01772_));
 sky130_vsdinv _20308_ (.A(net60),
    .Y(_01773_));
 sky130_vsdinv _20309_ (.A(net37),
    .Y(_01878_));
 sky130_fd_sc_hd__nand3b_1 _20310_ (.A_N(_14268_),
    .B(_15186_),
    .C(net46),
    .Y(_04106_));
 sky130_fd_sc_hd__nand3_1 _20311_ (.A(_15172_),
    .B(_14829_),
    .C(net54),
    .Y(_04107_));
 sky130_fd_sc_hd__o311a_1 _20312_ (.A1(_15169_),
    .A2(_15171_),
    .A3(_01878_),
    .B1(_04106_),
    .C1(_04107_),
    .X(_01774_));
 sky130_fd_sc_hd__o2bb2a_1 _20313_ (.A1_N(_04098_),
    .A2_N(_01776_),
    .B1(_01775_),
    .B2(_15201_),
    .X(_01777_));
 sky130_fd_sc_hd__and2_1 _20314_ (.A(_14185_),
    .B(_13679_),
    .X(_04108_));
 sky130_fd_sc_hd__a221oi_2 _20315_ (.A1(\count_instr[37] ),
    .A2(_14171_),
    .B1(\count_instr[5] ),
    .B2(_14183_),
    .C1(_04108_),
    .Y(_01781_));
 sky130_fd_sc_hd__and2_1 _20316_ (.A(_04085_),
    .B(\timer[5] ),
    .X(_04109_));
 sky130_fd_sc_hd__a221oi_2 _20317_ (.A1(\irq_mask[5] ),
    .A2(_14155_),
    .B1(\cpuregs_rs1[5] ),
    .B2(_15191_),
    .C1(_04109_),
    .Y(_01783_));
 sky130_fd_sc_hd__and2_1 _20318_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .X(_04110_));
 sky130_fd_sc_hd__nor2_4 _20319_ (.A(_13241_),
    .B(\decoded_imm[5] ),
    .Y(_04111_));
 sky130_fd_sc_hd__and2_1 _20320_ (.A(_13244_),
    .B(\decoded_imm[4] ),
    .X(_04112_));
 sky130_fd_sc_hd__a21oi_2 _20321_ (.A1(_04103_),
    .A2(_04102_),
    .B1(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__o31a_1 _20322_ (.A1(_04110_),
    .A2(_04111_),
    .A3(_04113_),
    .B1(_12845_),
    .X(_04114_));
 sky130_fd_sc_hd__o21ai_2 _20323_ (.A1(_04110_),
    .A2(_04111_),
    .B1(_04113_),
    .Y(_04115_));
 sky130_fd_sc_hd__a22oi_4 _20324_ (.A1(_15167_),
    .A2(_01779_),
    .B1(_04114_),
    .B2(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__o221ai_2 _20325_ (.A1(_15184_),
    .A2(_01784_),
    .B1(_12660_),
    .B2(_01778_),
    .C1(_04116_),
    .Y(_01785_));
 sky130_vsdinv _20326_ (.A(net61),
    .Y(_01786_));
 sky130_vsdinv _20327_ (.A(net38),
    .Y(_01891_));
 sky130_fd_sc_hd__nand3b_1 _20328_ (.A_N(_14268_),
    .B(_15186_),
    .C(net47),
    .Y(_04117_));
 sky130_fd_sc_hd__nand3_1 _20329_ (.A(_15172_),
    .B(_14829_),
    .C(net497),
    .Y(_04118_));
 sky130_fd_sc_hd__o311a_1 _20330_ (.A1(_14265_),
    .A2(_15170_),
    .A3(_01891_),
    .B1(_04117_),
    .C1(_04118_),
    .X(_01787_));
 sky130_fd_sc_hd__o2bb2a_1 _20331_ (.A1_N(_04098_),
    .A2_N(_01789_),
    .B1(_01788_),
    .B2(_15201_),
    .X(_01790_));
 sky130_fd_sc_hd__and2_1 _20332_ (.A(\count_instr[38] ),
    .B(_14170_),
    .X(_04119_));
 sky130_fd_sc_hd__a221oi_2 _20333_ (.A1(\count_instr[6] ),
    .A2(_04099_),
    .B1(_14186_),
    .B2(\count_cycle[38] ),
    .C1(_04119_),
    .Y(_01794_));
 sky130_fd_sc_hd__and2_1 _20334_ (.A(\irq_mask[6] ),
    .B(_15203_),
    .X(_04120_));
 sky130_fd_sc_hd__a221oi_2 _20335_ (.A1(_14139_),
    .A2(\timer[6] ),
    .B1(\cpuregs_rs1[6] ),
    .B2(_15191_),
    .C1(_04120_),
    .Y(_01796_));
 sky130_fd_sc_hd__xnor2_4 _20336_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .Y(_04121_));
 sky130_fd_sc_hd__o21ba_1 _20337_ (.A1(_04111_),
    .A2(_04113_),
    .B1_N(_04110_),
    .X(_04122_));
 sky130_fd_sc_hd__nor2_4 _20338_ (.A(_04121_),
    .B(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__and2_1 _20339_ (.A(_04122_),
    .B(_04121_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_2 _20340_ (.A(_12885_),
    .X(_04125_));
 sky130_fd_sc_hd__nand2_1 _20341_ (.A(_04125_),
    .B(_01792_),
    .Y(_04126_));
 sky130_fd_sc_hd__o221a_1 _20342_ (.A1(_01791_),
    .A2(_12659_),
    .B1(_13872_),
    .B2(_01797_),
    .C1(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__o31ai_1 _20343_ (.A1(_12813_),
    .A2(_04123_),
    .A3(_04124_),
    .B1(_04127_),
    .Y(_01798_));
 sky130_vsdinv _20344_ (.A(net62),
    .Y(_01799_));
 sky130_fd_sc_hd__nand3_1 _20345_ (.A(_14828_),
    .B(_14829_),
    .C(net57),
    .Y(_04128_));
 sky130_vsdinv _20346_ (.A(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__a221oi_2 _20347_ (.A1(_15160_),
    .A2(net500),
    .B1(net48),
    .B2(_15162_),
    .C1(_04129_),
    .Y(_01800_));
 sky130_fd_sc_hd__o2bb2a_1 _20348_ (.A1_N(_04098_),
    .A2_N(_01802_),
    .B1(_01801_),
    .B2(_15201_),
    .X(_01803_));
 sky130_fd_sc_hd__clkbuf_2 _20349_ (.A(instr_rdcycleh),
    .X(_04130_));
 sky130_fd_sc_hd__and2_1 _20350_ (.A(_04130_),
    .B(_13623_),
    .X(_04131_));
 sky130_fd_sc_hd__a221oi_2 _20351_ (.A1(\count_instr[39] ),
    .A2(_14171_),
    .B1(\count_instr[7] ),
    .B2(_14183_),
    .C1(_04131_),
    .Y(_01807_));
 sky130_fd_sc_hd__clkbuf_4 _20352_ (.A(_15190_),
    .X(_04132_));
 sky130_fd_sc_hd__and2_1 _20353_ (.A(_04085_),
    .B(\timer[7] ),
    .X(_04133_));
 sky130_fd_sc_hd__a221oi_2 _20354_ (.A1(\irq_mask[7] ),
    .A2(_14155_),
    .B1(\cpuregs_rs1[7] ),
    .B2(_04132_),
    .C1(_04133_),
    .Y(_01809_));
 sky130_fd_sc_hd__and2_2 _20355_ (.A(_13237_),
    .B(_14563_),
    .X(_04134_));
 sky130_fd_sc_hd__nor2_1 _20356_ (.A(\reg_pc[7] ),
    .B(_14566_),
    .Y(_04135_));
 sky130_fd_sc_hd__and2_1 _20357_ (.A(\reg_pc[7] ),
    .B(_14566_),
    .X(_04136_));
 sky130_fd_sc_hd__nor2_2 _20358_ (.A(_04135_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__o31a_1 _20359_ (.A1(_04134_),
    .A2(_04137_),
    .A3(_04123_),
    .B1(_14717_),
    .X(_04138_));
 sky130_fd_sc_hd__o21ai_1 _20360_ (.A1(_04134_),
    .A2(_04123_),
    .B1(_04137_),
    .Y(_04139_));
 sky130_vsdinv _20361_ (.A(_01804_),
    .Y(_04140_));
 sky130_fd_sc_hd__buf_4 _20362_ (.A(_12853_),
    .X(_04141_));
 sky130_fd_sc_hd__o2bb2ai_2 _20363_ (.A1_N(_12652_),
    .A2_N(_04140_),
    .B1(_01810_),
    .B2(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__a221o_1 _20364_ (.A1(_14827_),
    .A2(_01805_),
    .B1(_04138_),
    .B2(_04139_),
    .C1(_04142_),
    .X(_01811_));
 sky130_fd_sc_hd__clkbuf_2 _20365_ (.A(_15175_),
    .X(_04143_));
 sky130_fd_sc_hd__nand2_1 _20366_ (.A(_04143_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_4 _20367_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .Y(_01816_));
 sky130_vsdinv _20368_ (.A(latched_is_lh),
    .Y(_04144_));
 sky130_fd_sc_hd__clkbuf_2 _20369_ (.A(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__nand2_2 _20370_ (.A(_04140_),
    .B(latched_is_lb),
    .Y(_04146_));
 sky130_fd_sc_hd__clkbuf_2 _20371_ (.A(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__o21a_1 _20372_ (.A1(_04145_),
    .A2(_01815_),
    .B1(_04147_),
    .X(_01817_));
 sky130_fd_sc_hd__clkbuf_4 _20373_ (.A(_14185_),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_2 _20374_ (.A(instr_rdinstr),
    .X(_04149_));
 sky130_fd_sc_hd__and2_1 _20375_ (.A(\count_instr[8] ),
    .B(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__a221oi_2 _20376_ (.A1(\count_instr[40] ),
    .A2(_14171_),
    .B1(_04148_),
    .B2(_13599_),
    .C1(_04150_),
    .Y(_01821_));
 sky130_fd_sc_hd__clkbuf_4 _20377_ (.A(_12955_),
    .X(_04151_));
 sky130_fd_sc_hd__and2_1 _20378_ (.A(_04085_),
    .B(\timer[8] ),
    .X(_04152_));
 sky130_fd_sc_hd__a221oi_2 _20379_ (.A1(\irq_mask[8] ),
    .A2(_04151_),
    .B1(\cpuregs_rs1[8] ),
    .B2(_04132_),
    .C1(_04152_),
    .Y(_01823_));
 sky130_fd_sc_hd__xor2_4 _20380_ (.A(\reg_pc[8] ),
    .B(_14569_),
    .X(_04153_));
 sky130_fd_sc_hd__o21bai_1 _20381_ (.A1(_04134_),
    .A2(_04123_),
    .B1_N(_04135_),
    .Y(_04154_));
 sky130_fd_sc_hd__or2b_4 _20382_ (.A(_04136_),
    .B_N(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__xnor2_4 _20383_ (.A(_04153_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__a2bb2oi_4 _20384_ (.A1_N(_01824_),
    .A2_N(_04094_),
    .B1(_04080_),
    .B2(_01819_),
    .Y(_04157_));
 sky130_fd_sc_hd__o221ai_4 _20385_ (.A1(_04073_),
    .A2(_01818_),
    .B1(_12812_),
    .B2(_04156_),
    .C1(_04157_),
    .Y(_01825_));
 sky130_fd_sc_hd__nand2_1 _20386_ (.A(_04143_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__o21a_1 _20387_ (.A1(_04145_),
    .A2(_01829_),
    .B1(_04147_),
    .X(_01830_));
 sky130_fd_sc_hd__and2_1 _20388_ (.A(_04130_),
    .B(\count_cycle[41] ),
    .X(_04158_));
 sky130_fd_sc_hd__a221oi_2 _20389_ (.A1(\count_instr[41] ),
    .A2(_14171_),
    .B1(\count_instr[9] ),
    .B2(_14183_),
    .C1(_04158_),
    .Y(_01834_));
 sky130_fd_sc_hd__and2_1 _20390_ (.A(\irq_mask[9] ),
    .B(_15203_),
    .X(_04159_));
 sky130_fd_sc_hd__a221oi_2 _20391_ (.A1(_14139_),
    .A2(\timer[9] ),
    .B1(\cpuregs_rs1[9] ),
    .B2(_04132_),
    .C1(_04159_),
    .Y(_01836_));
 sky130_fd_sc_hd__and2_1 _20392_ (.A(\reg_pc[9] ),
    .B(_14571_),
    .X(_04160_));
 sky130_fd_sc_hd__nor2_2 _20393_ (.A(\reg_pc[9] ),
    .B(_14571_),
    .Y(_04161_));
 sky130_fd_sc_hd__and2_1 _20394_ (.A(\reg_pc[8] ),
    .B(_14569_),
    .X(_04162_));
 sky130_fd_sc_hd__a21oi_4 _20395_ (.A1(_04155_),
    .A2(_04153_),
    .B1(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__o31a_1 _20396_ (.A1(_04160_),
    .A2(_04161_),
    .A3(_04163_),
    .B1(_12845_),
    .X(_04164_));
 sky130_fd_sc_hd__o21ai_2 _20397_ (.A1(_04160_),
    .A2(_04161_),
    .B1(_04163_),
    .Y(_04165_));
 sky130_fd_sc_hd__a22oi_4 _20398_ (.A1(_15167_),
    .A2(_01832_),
    .B1(_04164_),
    .B2(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__o221ai_4 _20399_ (.A1(_15184_),
    .A2(_01837_),
    .B1(_12660_),
    .B2(_01831_),
    .C1(_04166_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_1 _20400_ (.A(_04143_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o21a_1 _20401_ (.A1(_04145_),
    .A2(_01842_),
    .B1(_04147_),
    .X(_01843_));
 sky130_fd_sc_hd__clkbuf_2 _20402_ (.A(instr_rdinstrh),
    .X(_04167_));
 sky130_fd_sc_hd__and2_1 _20403_ (.A(\count_instr[42] ),
    .B(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__a221oi_2 _20404_ (.A1(\count_instr[10] ),
    .A2(_04099_),
    .B1(_04148_),
    .B2(\count_cycle[42] ),
    .C1(_04168_),
    .Y(_01847_));
 sky130_fd_sc_hd__and2_1 _20405_ (.A(_04085_),
    .B(\timer[10] ),
    .X(_04169_));
 sky130_fd_sc_hd__a221oi_2 _20406_ (.A1(\irq_mask[10] ),
    .A2(_04151_),
    .B1(\cpuregs_rs1[10] ),
    .B2(_04132_),
    .C1(_04169_),
    .Y(_01849_));
 sky130_fd_sc_hd__and2_1 _20407_ (.A(\reg_pc[10] ),
    .B(\decoded_imm[10] ),
    .X(_04170_));
 sky130_fd_sc_hd__nor2_2 _20408_ (.A(\reg_pc[10] ),
    .B(\decoded_imm[10] ),
    .Y(_04171_));
 sky130_fd_sc_hd__o21ba_1 _20409_ (.A1(_04161_),
    .A2(_04163_),
    .B1_N(_04160_),
    .X(_04172_));
 sky130_fd_sc_hd__o21a_1 _20410_ (.A1(_04170_),
    .A2(_04171_),
    .B1(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__nor3_2 _20411_ (.A(_04170_),
    .B(_04171_),
    .C(_04172_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand2_1 _20412_ (.A(_04125_),
    .B(_01845_),
    .Y(_04175_));
 sky130_fd_sc_hd__o221a_2 _20413_ (.A1(_01844_),
    .A2(_12659_),
    .B1(_13872_),
    .B2(_01850_),
    .C1(_04175_),
    .X(_04176_));
 sky130_fd_sc_hd__o31ai_1 _20414_ (.A1(_15182_),
    .A2(_04173_),
    .A3(_04174_),
    .B1(_04176_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_1 _20415_ (.A(_04143_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__o21a_1 _20416_ (.A1(_04145_),
    .A2(_01855_),
    .B1(_04147_),
    .X(_01856_));
 sky130_fd_sc_hd__clkbuf_4 _20417_ (.A(instr_rdinstrh),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_4 _20418_ (.A(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__and2_1 _20419_ (.A(\count_instr[11] ),
    .B(_04149_),
    .X(_04179_));
 sky130_fd_sc_hd__a221oi_2 _20420_ (.A1(\count_instr[43] ),
    .A2(_04178_),
    .B1(_04148_),
    .B2(_13669_),
    .C1(_04179_),
    .Y(_01860_));
 sky130_fd_sc_hd__buf_1 _20421_ (.A(net494),
    .X(_04180_));
 sky130_fd_sc_hd__and2_1 _20422_ (.A(_04180_),
    .B(\timer[11] ),
    .X(_04181_));
 sky130_fd_sc_hd__a221oi_2 _20423_ (.A1(\irq_mask[11] ),
    .A2(_04151_),
    .B1(\cpuregs_rs1[11] ),
    .B2(_04132_),
    .C1(_04181_),
    .Y(_01862_));
 sky130_fd_sc_hd__o21ba_1 _20424_ (.A1(_04171_),
    .A2(_04172_),
    .B1_N(_04170_),
    .X(_04182_));
 sky130_fd_sc_hd__xnor2_4 _20425_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .Y(_04183_));
 sky130_fd_sc_hd__and2_1 _20426_ (.A(_04182_),
    .B(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__o21bai_2 _20427_ (.A1(_04183_),
    .A2(_04182_),
    .B1_N(_12811_),
    .Y(_04185_));
 sky130_fd_sc_hd__a2bb2oi_4 _20428_ (.A1_N(_01863_),
    .A2_N(_04094_),
    .B1(_04080_),
    .B2(_01858_),
    .Y(_04186_));
 sky130_fd_sc_hd__o221ai_4 _20429_ (.A1(_04073_),
    .A2(_01857_),
    .B1(_04184_),
    .B2(_04185_),
    .C1(_04186_),
    .Y(_01864_));
 sky130_fd_sc_hd__nand2_1 _20430_ (.A(_04143_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__o21a_1 _20431_ (.A1(_04145_),
    .A2(_01868_),
    .B1(_04147_),
    .X(_01869_));
 sky130_fd_sc_hd__and2_1 _20432_ (.A(_04130_),
    .B(\count_cycle[44] ),
    .X(_04187_));
 sky130_fd_sc_hd__a221oi_2 _20433_ (.A1(\count_instr[44] ),
    .A2(_04178_),
    .B1(\count_instr[12] ),
    .B2(_14183_),
    .C1(_04187_),
    .Y(_01873_));
 sky130_fd_sc_hd__and2_1 _20434_ (.A(\irq_mask[12] ),
    .B(_15203_),
    .X(_04188_));
 sky130_fd_sc_hd__a221oi_2 _20435_ (.A1(_14139_),
    .A2(\timer[12] ),
    .B1(\cpuregs_rs1[12] ),
    .B2(_04132_),
    .C1(_04188_),
    .Y(_01875_));
 sky130_fd_sc_hd__and2_1 _20436_ (.A(\reg_pc[12] ),
    .B(\decoded_imm[12] ),
    .X(_04189_));
 sky130_fd_sc_hd__nor2_2 _20437_ (.A(\reg_pc[12] ),
    .B(\decoded_imm[12] ),
    .Y(_04190_));
 sky130_fd_sc_hd__and2_1 _20438_ (.A(_13223_),
    .B(\decoded_imm[11] ),
    .X(_04191_));
 sky130_fd_sc_hd__o21ba_1 _20439_ (.A1(_04183_),
    .A2(_04182_),
    .B1_N(_04191_),
    .X(_04192_));
 sky130_fd_sc_hd__o21a_1 _20440_ (.A1(_04189_),
    .A2(_04190_),
    .B1(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__nor3_2 _20441_ (.A(_04189_),
    .B(_04190_),
    .C(_04192_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _20442_ (.A(_12843_),
    .B(_01871_),
    .Y(_04195_));
 sky130_fd_sc_hd__o221a_2 _20443_ (.A1(_01870_),
    .A2(_12659_),
    .B1(_13872_),
    .B2(_01876_),
    .C1(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__o31ai_1 _20444_ (.A1(_15182_),
    .A2(_04193_),
    .A3(_04194_),
    .B1(_04196_),
    .Y(_01877_));
 sky130_fd_sc_hd__nand2_1 _20445_ (.A(_04143_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__o21a_1 _20446_ (.A1(_04145_),
    .A2(_01881_),
    .B1(_04147_),
    .X(_01882_));
 sky130_fd_sc_hd__and2_1 _20447_ (.A(\count_instr[13] ),
    .B(_04149_),
    .X(_04197_));
 sky130_fd_sc_hd__a221oi_2 _20448_ (.A1(\count_instr[45] ),
    .A2(_04178_),
    .B1(_04148_),
    .B2(_13626_),
    .C1(_04197_),
    .Y(_01886_));
 sky130_fd_sc_hd__clkbuf_4 _20449_ (.A(_15190_),
    .X(_04198_));
 sky130_fd_sc_hd__and2_1 _20450_ (.A(_04180_),
    .B(\timer[13] ),
    .X(_04199_));
 sky130_fd_sc_hd__a221oi_2 _20451_ (.A1(\irq_mask[13] ),
    .A2(_04151_),
    .B1(\cpuregs_rs1[13] ),
    .B2(_04198_),
    .C1(_04199_),
    .Y(_01888_));
 sky130_fd_sc_hd__and2_1 _20452_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .X(_04200_));
 sky130_vsdinv _20453_ (.A(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__or2_2 _20454_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .X(_04202_));
 sky130_fd_sc_hd__o21bai_2 _20455_ (.A1(_04190_),
    .A2(_04192_),
    .B1_N(_04189_),
    .Y(_04203_));
 sky130_fd_sc_hd__a21o_1 _20456_ (.A1(_04201_),
    .A2(_04202_),
    .B1(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__nand3_1 _20457_ (.A(_04203_),
    .B(_04201_),
    .C(_04202_),
    .Y(_04205_));
 sky130_fd_sc_hd__and2b_1 _20458_ (.A_N(_01883_),
    .B(_13092_),
    .X(_04206_));
 sky130_fd_sc_hd__o2bb2ai_4 _20459_ (.A1_N(_14713_),
    .A2_N(_01884_),
    .B1(_01889_),
    .B2(_04141_),
    .Y(_04207_));
 sky130_fd_sc_hd__a311o_1 _20460_ (.A1(_04204_),
    .A2(_04205_),
    .A3(_14718_),
    .B1(_04206_),
    .C1(_04207_),
    .X(_01890_));
 sky130_fd_sc_hd__nand2_1 _20461_ (.A(_15176_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__o21a_1 _20462_ (.A1(_04144_),
    .A2(_01894_),
    .B1(_04146_),
    .X(_01895_));
 sky130_vsdinv _20463_ (.A(\count_cycle[14] ),
    .Y(_01898_));
 sky130_fd_sc_hd__and2_1 _20464_ (.A(\count_instr[46] ),
    .B(_04167_),
    .X(_04208_));
 sky130_fd_sc_hd__a221oi_2 _20465_ (.A1(\count_instr[14] ),
    .A2(_04099_),
    .B1(_04148_),
    .B2(_13602_),
    .C1(_04208_),
    .Y(_01899_));
 sky130_fd_sc_hd__clkbuf_4 _20466_ (.A(_14138_),
    .X(_04209_));
 sky130_fd_sc_hd__and2_1 _20467_ (.A(\irq_mask[14] ),
    .B(_15203_),
    .X(_04210_));
 sky130_fd_sc_hd__a221oi_2 _20468_ (.A1(_04209_),
    .A2(\timer[14] ),
    .B1(\cpuregs_rs1[14] ),
    .B2(_04198_),
    .C1(_04210_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_2 _20469_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .Y(_04211_));
 sky130_fd_sc_hd__and2_1 _20470_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .X(_04212_));
 sky130_fd_sc_hd__nor2_2 _20471_ (.A(_04211_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__a21oi_4 _20472_ (.A1(_04203_),
    .A2(_04202_),
    .B1(_04200_),
    .Y(_04214_));
 sky130_fd_sc_hd__xor2_2 _20473_ (.A(_04213_),
    .B(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_4 _20474_ (.A(_12658_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_4 _20475_ (.A(_12853_),
    .X(_04217_));
 sky130_fd_sc_hd__nand2_1 _20476_ (.A(_04125_),
    .B(_01897_),
    .Y(_04218_));
 sky130_fd_sc_hd__o221ai_4 _20477_ (.A1(_01896_),
    .A2(_04216_),
    .B1(_01902_),
    .B2(_04217_),
    .C1(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__o21bai_1 _20478_ (.A1(_12813_),
    .A2(_04215_),
    .B1_N(_04219_),
    .Y(_01903_));
 sky130_vsdinv _20479_ (.A(net500),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_1 _20480_ (.A(_15176_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__o21a_4 _20481_ (.A1(_04144_),
    .A2(_01907_),
    .B1(_04146_),
    .X(_01908_));
 sky130_vsdinv _20482_ (.A(\count_cycle[15] ),
    .Y(_01911_));
 sky130_fd_sc_hd__and2_1 _20483_ (.A(\count_instr[15] ),
    .B(_04149_),
    .X(_04220_));
 sky130_fd_sc_hd__a221oi_2 _20484_ (.A1(\count_instr[47] ),
    .A2(_04178_),
    .B1(_04148_),
    .B2(\count_cycle[47] ),
    .C1(_04220_),
    .Y(_01912_));
 sky130_fd_sc_hd__and2_1 _20485_ (.A(\irq_mask[15] ),
    .B(_15203_),
    .X(_04221_));
 sky130_fd_sc_hd__a221oi_2 _20486_ (.A1(_04209_),
    .A2(\timer[15] ),
    .B1(\cpuregs_rs1[15] ),
    .B2(_04198_),
    .C1(_04221_),
    .Y(_01914_));
 sky130_fd_sc_hd__and2_1 _20487_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .X(_04222_));
 sky130_vsdinv _20488_ (.A(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__or2_2 _20489_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .X(_04224_));
 sky130_fd_sc_hd__o21bai_2 _20490_ (.A1(_04211_),
    .A2(_04214_),
    .B1_N(_04212_),
    .Y(_04225_));
 sky130_fd_sc_hd__a21o_1 _20491_ (.A1(_04223_),
    .A2(_04224_),
    .B1(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__nand3_4 _20492_ (.A(_04225_),
    .B(_04223_),
    .C(_04224_),
    .Y(_04227_));
 sky130_fd_sc_hd__and2b_1 _20493_ (.A_N(_01909_),
    .B(_13092_),
    .X(_04228_));
 sky130_fd_sc_hd__o2bb2ai_4 _20494_ (.A1_N(_14713_),
    .A2_N(_01910_),
    .B1(_01915_),
    .B2(_04141_),
    .Y(_04229_));
 sky130_fd_sc_hd__a311o_1 _20495_ (.A1(_04226_),
    .A2(_04227_),
    .A3(_14718_),
    .B1(_04228_),
    .C1(_04229_),
    .X(_01916_));
 sky130_fd_sc_hd__clkbuf_2 _20496_ (.A(_14818_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_2 _20497_ (.A(_14833_),
    .X(_04231_));
 sky130_fd_sc_hd__nand3_1 _20498_ (.A(_04230_),
    .B(_04231_),
    .C(net40),
    .Y(_01917_));
 sky130_vsdinv _20499_ (.A(_13613_),
    .Y(_01920_));
 sky130_fd_sc_hd__clkbuf_4 _20500_ (.A(_14182_),
    .X(_04232_));
 sky130_fd_sc_hd__and2_1 _20501_ (.A(_04130_),
    .B(_13628_),
    .X(_04233_));
 sky130_fd_sc_hd__a221oi_2 _20502_ (.A1(\count_instr[48] ),
    .A2(_04178_),
    .B1(\count_instr[16] ),
    .B2(_04232_),
    .C1(_04233_),
    .Y(_01921_));
 sky130_fd_sc_hd__and2_1 _20503_ (.A(_04180_),
    .B(\timer[16] ),
    .X(_04234_));
 sky130_fd_sc_hd__a221oi_2 _20504_ (.A1(\irq_mask[16] ),
    .A2(_04151_),
    .B1(\cpuregs_rs1[16] ),
    .B2(_04198_),
    .C1(_04234_),
    .Y(_01923_));
 sky130_fd_sc_hd__xor2_4 _20505_ (.A(\reg_pc[16] ),
    .B(\decoded_imm[16] ),
    .X(_04235_));
 sky130_fd_sc_hd__a21bo_1 _20506_ (.A1(_04227_),
    .A2(_04223_),
    .B1_N(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__nand3b_1 _20507_ (.A_N(_04235_),
    .B(_04227_),
    .C(_04223_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_2 _20508_ (.A(_04125_),
    .B(_01919_),
    .Y(_04238_));
 sky130_fd_sc_hd__o221ai_4 _20509_ (.A1(_01918_),
    .A2(_04216_),
    .B1(_01924_),
    .B2(_04141_),
    .C1(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__a31o_1 _20510_ (.A1(_04236_),
    .A2(_14822_),
    .A3(_04237_),
    .B1(_04239_),
    .X(_01925_));
 sky130_fd_sc_hd__nand3_1 _20511_ (.A(_04230_),
    .B(_04231_),
    .C(net499),
    .Y(_01926_));
 sky130_vsdinv _20512_ (.A(\count_cycle[17] ),
    .Y(_01929_));
 sky130_fd_sc_hd__clkbuf_4 _20513_ (.A(_14185_),
    .X(_04240_));
 sky130_fd_sc_hd__and2_1 _20514_ (.A(\count_instr[49] ),
    .B(_04167_),
    .X(_04241_));
 sky130_fd_sc_hd__a221oi_2 _20515_ (.A1(\count_instr[17] ),
    .A2(_04099_),
    .B1(_04240_),
    .B2(_13661_),
    .C1(_04241_),
    .Y(_01930_));
 sky130_fd_sc_hd__and2_1 _20516_ (.A(_04180_),
    .B(\timer[17] ),
    .X(_04242_));
 sky130_fd_sc_hd__a221oi_2 _20517_ (.A1(\irq_mask[17] ),
    .A2(_04151_),
    .B1(\cpuregs_rs1[17] ),
    .B2(_04198_),
    .C1(_04242_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_2 _20518_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .Y(_04243_));
 sky130_fd_sc_hd__and2_2 _20519_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .X(_04244_));
 sky130_fd_sc_hd__nor2_4 _20520_ (.A(_04243_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__and2_1 _20521_ (.A(_13205_),
    .B(_14594_),
    .X(_04246_));
 sky130_fd_sc_hd__or2b_1 _20522_ (.A(_04246_),
    .B_N(_04236_),
    .X(_04247_));
 sky130_fd_sc_hd__o21a_1 _20523_ (.A1(_04245_),
    .A2(_04247_),
    .B1(_14717_),
    .X(_04248_));
 sky130_fd_sc_hd__nand2_1 _20524_ (.A(_04247_),
    .B(_04245_),
    .Y(_04249_));
 sky130_fd_sc_hd__a22oi_4 _20525_ (.A1(_15167_),
    .A2(_01928_),
    .B1(_04248_),
    .B2(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__o221ai_4 _20526_ (.A1(_15184_),
    .A2(_01933_),
    .B1(_12660_),
    .B2(_01927_),
    .C1(_04250_),
    .Y(_01934_));
 sky130_fd_sc_hd__nand3_1 _20527_ (.A(_04230_),
    .B(_04231_),
    .C(net42),
    .Y(_01935_));
 sky130_vsdinv _20528_ (.A(\count_cycle[18] ),
    .Y(_01938_));
 sky130_fd_sc_hd__and2_1 _20529_ (.A(\count_instr[50] ),
    .B(_04167_),
    .X(_04251_));
 sky130_fd_sc_hd__a221oi_2 _20530_ (.A1(\count_instr[18] ),
    .A2(_04099_),
    .B1(_04240_),
    .B2(_13604_),
    .C1(_04251_),
    .Y(_01939_));
 sky130_fd_sc_hd__buf_1 _20531_ (.A(_12908_),
    .X(_04252_));
 sky130_fd_sc_hd__and2_1 _20532_ (.A(\irq_mask[18] ),
    .B(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__a221oi_2 _20533_ (.A1(_04209_),
    .A2(\timer[18] ),
    .B1(\cpuregs_rs1[18] ),
    .B2(_04198_),
    .C1(_04253_),
    .Y(_01941_));
 sky130_fd_sc_hd__nand2_1 _20534_ (.A(_04235_),
    .B(_04245_),
    .Y(_04254_));
 sky130_fd_sc_hd__a21o_1 _20535_ (.A1(_04227_),
    .A2(_04223_),
    .B1(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__o211a_1 _20536_ (.A1(\reg_pc[17] ),
    .A2(_14597_),
    .B1(\reg_pc[16] ),
    .C1(_14594_),
    .X(_04256_));
 sky130_fd_sc_hd__nor2_4 _20537_ (.A(_04244_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__xnor2_1 _20538_ (.A(_13199_),
    .B(_14600_),
    .Y(_04258_));
 sky130_fd_sc_hd__a21o_1 _20539_ (.A1(_04255_),
    .A2(_04257_),
    .B1(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__nand3_1 _20540_ (.A(_04255_),
    .B(_04258_),
    .C(_04257_),
    .Y(_04260_));
 sky130_fd_sc_hd__and2b_1 _20541_ (.A_N(_01936_),
    .B(_13092_),
    .X(_04261_));
 sky130_fd_sc_hd__o2bb2ai_4 _20542_ (.A1_N(_14713_),
    .A2_N(_01937_),
    .B1(_01942_),
    .B2(_04141_),
    .Y(_04262_));
 sky130_fd_sc_hd__a311o_1 _20543_ (.A1(_04259_),
    .A2(_14718_),
    .A3(_04260_),
    .B1(_04261_),
    .C1(_04262_),
    .X(_01943_));
 sky130_fd_sc_hd__nand3_1 _20544_ (.A(_04230_),
    .B(_04231_),
    .C(net498),
    .Y(_01944_));
 sky130_vsdinv _20545_ (.A(_13588_),
    .Y(_01947_));
 sky130_fd_sc_hd__and2_1 _20546_ (.A(_04130_),
    .B(_13656_),
    .X(_04263_));
 sky130_fd_sc_hd__a221oi_2 _20547_ (.A1(\count_instr[51] ),
    .A2(_04178_),
    .B1(\count_instr[19] ),
    .B2(_04232_),
    .C1(_04263_),
    .Y(_01948_));
 sky130_fd_sc_hd__clkbuf_4 _20548_ (.A(_12955_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_4 _20549_ (.A(_15190_),
    .X(_04265_));
 sky130_fd_sc_hd__and2_1 _20550_ (.A(_04180_),
    .B(\timer[19] ),
    .X(_04266_));
 sky130_fd_sc_hd__a221oi_2 _20551_ (.A1(\irq_mask[19] ),
    .A2(_04264_),
    .B1(\cpuregs_rs1[19] ),
    .B2(_04265_),
    .C1(_04266_),
    .Y(_01950_));
 sky130_vsdinv _20552_ (.A(\reg_pc[18] ),
    .Y(_04267_));
 sky130_vsdinv _20553_ (.A(\decoded_imm[18] ),
    .Y(_04268_));
 sky130_fd_sc_hd__and2_1 _20554_ (.A(\reg_pc[19] ),
    .B(\decoded_imm[19] ),
    .X(_04269_));
 sky130_fd_sc_hd__nor2_8 _20555_ (.A(\reg_pc[19] ),
    .B(\decoded_imm[19] ),
    .Y(_04270_));
 sky130_fd_sc_hd__o221a_1 _20556_ (.A1(_04267_),
    .A2(_04268_),
    .B1(_04269_),
    .B2(_04270_),
    .C1(_04259_),
    .X(_04271_));
 sky130_fd_sc_hd__nand2_1 _20557_ (.A(_04255_),
    .B(_04257_),
    .Y(_04272_));
 sky130_fd_sc_hd__nand2_1 _20558_ (.A(_04267_),
    .B(_04268_),
    .Y(_04273_));
 sky130_fd_sc_hd__and2_1 _20559_ (.A(\reg_pc[18] ),
    .B(_14600_),
    .X(_04274_));
 sky130_fd_sc_hd__a21oi_4 _20560_ (.A1(_04272_),
    .A2(_04273_),
    .B1(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__o31ai_4 _20561_ (.A1(_04269_),
    .A2(_04270_),
    .A3(_04275_),
    .B1(_04092_),
    .Y(_04276_));
 sky130_fd_sc_hd__a2bb2oi_4 _20562_ (.A1_N(_01951_),
    .A2_N(_04094_),
    .B1(_04080_),
    .B2(_01946_),
    .Y(_04277_));
 sky130_fd_sc_hd__o221ai_4 _20563_ (.A1(_04073_),
    .A2(_01945_),
    .B1(_04271_),
    .B2(_04276_),
    .C1(_04277_),
    .Y(_01952_));
 sky130_fd_sc_hd__nand3_1 _20564_ (.A(_04230_),
    .B(_04231_),
    .C(net45),
    .Y(_01953_));
 sky130_vsdinv _20565_ (.A(\count_cycle[20] ),
    .Y(_01956_));
 sky130_fd_sc_hd__clkbuf_4 _20566_ (.A(_04177_),
    .X(_04278_));
 sky130_fd_sc_hd__and2_1 _20567_ (.A(\count_instr[20] ),
    .B(_04149_),
    .X(_04279_));
 sky130_fd_sc_hd__a221oi_2 _20568_ (.A1(\count_instr[52] ),
    .A2(_04278_),
    .B1(_04240_),
    .B2(_13654_),
    .C1(_04279_),
    .Y(_01957_));
 sky130_fd_sc_hd__and2_1 _20569_ (.A(\irq_mask[20] ),
    .B(_04252_),
    .X(_04280_));
 sky130_fd_sc_hd__a221oi_2 _20570_ (.A1(_04209_),
    .A2(\timer[20] ),
    .B1(\cpuregs_rs1[20] ),
    .B2(_04265_),
    .C1(_04280_),
    .Y(_01959_));
 sky130_fd_sc_hd__a2bb2oi_4 _20571_ (.A1_N(_01960_),
    .A2_N(_15197_),
    .B1(_13548_),
    .B2(_01955_),
    .Y(_04281_));
 sky130_fd_sc_hd__and2_1 _20572_ (.A(\reg_pc[20] ),
    .B(\decoded_imm[20] ),
    .X(_04282_));
 sky130_vsdinv _20573_ (.A(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__or2_2 _20574_ (.A(\reg_pc[20] ),
    .B(\decoded_imm[20] ),
    .X(_04284_));
 sky130_fd_sc_hd__o21bai_4 _20575_ (.A1(_04270_),
    .A2(_04275_),
    .B1_N(_04269_),
    .Y(_04285_));
 sky130_fd_sc_hd__a21o_1 _20576_ (.A1(_04283_),
    .A2(_04284_),
    .B1(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__nand3_2 _20577_ (.A(_04285_),
    .B(_04283_),
    .C(_04284_),
    .Y(_04287_));
 sky130_fd_sc_hd__nand3_4 _20578_ (.A(_04286_),
    .B(_04092_),
    .C(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__o211ai_4 _20579_ (.A1(_15181_),
    .A2(_01954_),
    .B1(_04281_),
    .C1(_04288_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand3_1 _20580_ (.A(_04230_),
    .B(_04231_),
    .C(net46),
    .Y(_01962_));
 sky130_vsdinv _20581_ (.A(\count_cycle[21] ),
    .Y(_01965_));
 sky130_fd_sc_hd__and2_1 _20582_ (.A(_04130_),
    .B(\count_cycle[53] ),
    .X(_04289_));
 sky130_fd_sc_hd__a221oi_2 _20583_ (.A1(\count_instr[53] ),
    .A2(_04278_),
    .B1(\count_instr[21] ),
    .B2(_04232_),
    .C1(_04289_),
    .Y(_01966_));
 sky130_fd_sc_hd__and2_1 _20584_ (.A(_04180_),
    .B(\timer[21] ),
    .X(_04290_));
 sky130_fd_sc_hd__a221oi_2 _20585_ (.A1(\irq_mask[21] ),
    .A2(_04264_),
    .B1(\cpuregs_rs1[21] ),
    .B2(_04265_),
    .C1(_04290_),
    .Y(_01968_));
 sky130_fd_sc_hd__nor2_4 _20586_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .Y(_04291_));
 sky130_fd_sc_hd__and2_1 _20587_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .X(_04292_));
 sky130_fd_sc_hd__nor2_4 _20588_ (.A(_04291_),
    .B(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__a21oi_4 _20589_ (.A1(_04285_),
    .A2(_04284_),
    .B1(_04282_),
    .Y(_04294_));
 sky130_fd_sc_hd__xor2_4 _20590_ (.A(_04293_),
    .B(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__a2bb2oi_4 _20591_ (.A1_N(_01969_),
    .A2_N(_04094_),
    .B1(_13548_),
    .B2(_01964_),
    .Y(_04296_));
 sky130_fd_sc_hd__o221ai_4 _20592_ (.A1(_12660_),
    .A2(_01963_),
    .B1(_12812_),
    .B2(_04295_),
    .C1(_04296_),
    .Y(_01970_));
 sky130_fd_sc_hd__clkbuf_2 _20593_ (.A(_14817_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_2 _20594_ (.A(_14833_),
    .X(_04298_));
 sky130_fd_sc_hd__nand3_1 _20595_ (.A(_04297_),
    .B(_04298_),
    .C(net47),
    .Y(_01971_));
 sky130_vsdinv _20596_ (.A(_13590_),
    .Y(_01974_));
 sky130_fd_sc_hd__buf_1 _20597_ (.A(instr_rdcycleh),
    .X(_04299_));
 sky130_fd_sc_hd__and2_1 _20598_ (.A(_04299_),
    .B(\count_cycle[54] ),
    .X(_04300_));
 sky130_fd_sc_hd__a221oi_2 _20599_ (.A1(\count_instr[54] ),
    .A2(_04278_),
    .B1(\count_instr[22] ),
    .B2(_04232_),
    .C1(_04300_),
    .Y(_01975_));
 sky130_fd_sc_hd__and2_1 _20600_ (.A(_14137_),
    .B(\timer[22] ),
    .X(_04301_));
 sky130_fd_sc_hd__a221oi_2 _20601_ (.A1(\irq_mask[22] ),
    .A2(_04264_),
    .B1(\cpuregs_rs1[22] ),
    .B2(_04265_),
    .C1(_04301_),
    .Y(_01977_));
 sky130_fd_sc_hd__a2bb2oi_4 _20602_ (.A1_N(_01978_),
    .A2_N(_15197_),
    .B1(_13548_),
    .B2(_01973_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_4 _20603_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .Y(_04303_));
 sky130_fd_sc_hd__or2_2 _20604_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .X(_04304_));
 sky130_fd_sc_hd__o21bai_2 _20605_ (.A1(_04291_),
    .A2(_04294_),
    .B1_N(_04292_),
    .Y(_04305_));
 sky130_fd_sc_hd__a21o_1 _20606_ (.A1(_04303_),
    .A2(_04304_),
    .B1(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__nand3_4 _20607_ (.A(_04305_),
    .B(_04303_),
    .C(_04304_),
    .Y(_04307_));
 sky130_fd_sc_hd__nand3_4 _20608_ (.A(_04306_),
    .B(_04092_),
    .C(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__o211ai_4 _20609_ (.A1(_15181_),
    .A2(_01972_),
    .B1(_04302_),
    .C1(_04308_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand3_1 _20610_ (.A(_04297_),
    .B(_04298_),
    .C(net48),
    .Y(_01980_));
 sky130_vsdinv _20611_ (.A(\count_cycle[23] ),
    .Y(_01983_));
 sky130_fd_sc_hd__and2_1 _20612_ (.A(\count_instr[23] ),
    .B(_04149_),
    .X(_04309_));
 sky130_fd_sc_hd__a221oi_2 _20613_ (.A1(\count_instr[55] ),
    .A2(_04278_),
    .B1(_04240_),
    .B2(_13636_),
    .C1(_04309_),
    .Y(_01984_));
 sky130_fd_sc_hd__and2_1 _20614_ (.A(\irq_mask[23] ),
    .B(_04252_),
    .X(_04310_));
 sky130_fd_sc_hd__a221oi_2 _20615_ (.A1(_04209_),
    .A2(\timer[23] ),
    .B1(\cpuregs_rs1[23] ),
    .B2(_04265_),
    .C1(_04310_),
    .Y(_01986_));
 sky130_fd_sc_hd__a2bb2oi_4 _20616_ (.A1_N(_01987_),
    .A2_N(_15197_),
    .B1(_13548_),
    .B2(_01982_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand2_1 _20617_ (.A(_04307_),
    .B(_04303_),
    .Y(_04312_));
 sky130_fd_sc_hd__xor2_4 _20618_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .X(_04313_));
 sky130_fd_sc_hd__nand2_1 _20619_ (.A(_04312_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__nand3b_4 _20620_ (.A_N(_04313_),
    .B(_04307_),
    .C(_04303_),
    .Y(_04315_));
 sky130_fd_sc_hd__nand3_4 _20621_ (.A(_04314_),
    .B(_04092_),
    .C(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__o211ai_4 _20622_ (.A1(_15181_),
    .A2(_01981_),
    .B1(_04311_),
    .C1(_04316_),
    .Y(_01988_));
 sky130_fd_sc_hd__nand3_1 _20623_ (.A(_04297_),
    .B(_04298_),
    .C(net49),
    .Y(_01989_));
 sky130_vsdinv _20624_ (.A(_13617_),
    .Y(_01992_));
 sky130_fd_sc_hd__and2_1 _20625_ (.A(_04299_),
    .B(_13647_),
    .X(_04317_));
 sky130_fd_sc_hd__a221oi_2 _20626_ (.A1(\count_instr[56] ),
    .A2(_04278_),
    .B1(\count_instr[24] ),
    .B2(_04232_),
    .C1(_04317_),
    .Y(_01993_));
 sky130_fd_sc_hd__and2_1 _20627_ (.A(\irq_mask[24] ),
    .B(_04252_),
    .X(_04318_));
 sky130_fd_sc_hd__a221oi_2 _20628_ (.A1(_04209_),
    .A2(\timer[24] ),
    .B1(\cpuregs_rs1[24] ),
    .B2(_04265_),
    .C1(_04318_),
    .Y(_01995_));
 sky130_fd_sc_hd__and2_1 _20629_ (.A(_13182_),
    .B(\decoded_imm[23] ),
    .X(_04319_));
 sky130_fd_sc_hd__xor2_2 _20630_ (.A(\reg_pc[24] ),
    .B(_14615_),
    .X(_04320_));
 sky130_fd_sc_hd__a211o_1 _20631_ (.A1(_04312_),
    .A2(_04313_),
    .B1(_04319_),
    .C1(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__a21o_1 _20632_ (.A1(_04312_),
    .A2(_04313_),
    .B1(_04319_),
    .X(_04322_));
 sky130_fd_sc_hd__nand2_1 _20633_ (.A(_04322_),
    .B(_04320_),
    .Y(_04323_));
 sky130_fd_sc_hd__and2b_1 _20634_ (.A_N(_01990_),
    .B(_13092_),
    .X(_04324_));
 sky130_fd_sc_hd__o2bb2ai_2 _20635_ (.A1_N(_14713_),
    .A2_N(_01991_),
    .B1(_01996_),
    .B2(_04141_),
    .Y(_04325_));
 sky130_fd_sc_hd__a311o_2 _20636_ (.A1(_04321_),
    .A2(_04323_),
    .A3(_14718_),
    .B1(_04324_),
    .C1(_04325_),
    .X(_01997_));
 sky130_fd_sc_hd__nand3_1 _20637_ (.A(_04297_),
    .B(_04298_),
    .C(net50),
    .Y(_01998_));
 sky130_vsdinv _20638_ (.A(_13697_),
    .Y(_02001_));
 sky130_fd_sc_hd__and2_1 _20639_ (.A(_04299_),
    .B(_13638_),
    .X(_04326_));
 sky130_fd_sc_hd__a221oi_2 _20640_ (.A1(\count_instr[57] ),
    .A2(_04278_),
    .B1(\count_instr[25] ),
    .B2(_04232_),
    .C1(_04326_),
    .Y(_02002_));
 sky130_fd_sc_hd__clkbuf_4 _20641_ (.A(_15190_),
    .X(_04327_));
 sky130_fd_sc_hd__and2_1 _20642_ (.A(_14137_),
    .B(\timer[25] ),
    .X(_04328_));
 sky130_fd_sc_hd__a221oi_2 _20643_ (.A1(\irq_mask[25] ),
    .A2(_04264_),
    .B1(\cpuregs_rs1[25] ),
    .B2(_04327_),
    .C1(_04328_),
    .Y(_02004_));
 sky130_fd_sc_hd__and2_1 _20644_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .X(_04329_));
 sky130_vsdinv _20645_ (.A(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__nor2_1 _20646_ (.A(\reg_pc[25] ),
    .B(_14618_),
    .Y(_04331_));
 sky130_fd_sc_hd__and2_1 _20647_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .X(_04332_));
 sky130_fd_sc_hd__nor2_1 _20648_ (.A(_04331_),
    .B(_04332_),
    .Y(_04333_));
 sky130_vsdinv _20649_ (.A(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__a31oi_1 _20650_ (.A1(_04323_),
    .A2(_04330_),
    .A3(_04334_),
    .B1(_12812_),
    .Y(_04335_));
 sky130_fd_sc_hd__a21o_1 _20651_ (.A1(_04323_),
    .A2(_04330_),
    .B1(_04334_),
    .X(_04336_));
 sky130_fd_sc_hd__o22ai_2 _20652_ (.A1(_01999_),
    .A2(_04216_),
    .B1(_04217_),
    .B2(_02005_),
    .Y(_04337_));
 sky130_fd_sc_hd__a221o_2 _20653_ (.A1(_14827_),
    .A2(_02000_),
    .B1(_04335_),
    .B2(_04336_),
    .C1(_04337_),
    .X(_02006_));
 sky130_fd_sc_hd__nand3_1 _20654_ (.A(_04297_),
    .B(_04298_),
    .C(net51),
    .Y(_02007_));
 sky130_vsdinv _20655_ (.A(\count_cycle[26] ),
    .Y(_02010_));
 sky130_fd_sc_hd__and2_1 _20656_ (.A(_04299_),
    .B(_13642_),
    .X(_04338_));
 sky130_fd_sc_hd__a221oi_2 _20657_ (.A1(\count_instr[58] ),
    .A2(_04177_),
    .B1(\count_instr[26] ),
    .B2(_15178_),
    .C1(_04338_),
    .Y(_02011_));
 sky130_fd_sc_hd__and2_1 _20658_ (.A(\irq_mask[26] ),
    .B(_04252_),
    .X(_04339_));
 sky130_fd_sc_hd__a221oi_2 _20659_ (.A1(_14138_),
    .A2(\timer[26] ),
    .B1(\cpuregs_rs1[26] ),
    .B2(_04327_),
    .C1(_04339_),
    .Y(_02013_));
 sky130_fd_sc_hd__and2_1 _20660_ (.A(_04320_),
    .B(_04333_),
    .X(_04340_));
 sky130_fd_sc_hd__o21ba_1 _20661_ (.A1(_04331_),
    .A2(_04330_),
    .B1_N(_04332_),
    .X(_04341_));
 sky130_fd_sc_hd__a21boi_4 _20662_ (.A1(_04322_),
    .A2(_04340_),
    .B1_N(_04341_),
    .Y(_04342_));
 sky130_fd_sc_hd__xor2_2 _20663_ (.A(\reg_pc[26] ),
    .B(\decoded_imm[26] ),
    .X(_04343_));
 sky130_fd_sc_hd__or2b_1 _20664_ (.A(_04342_),
    .B_N(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__or2b_1 _20665_ (.A(_04343_),
    .B_N(_04342_),
    .X(_04345_));
 sky130_fd_sc_hd__nand2_1 _20666_ (.A(_04125_),
    .B(_02009_),
    .Y(_04346_));
 sky130_fd_sc_hd__o221ai_2 _20667_ (.A1(_02008_),
    .A2(_04216_),
    .B1(_02014_),
    .B2(_04217_),
    .C1(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__a31o_1 _20668_ (.A1(_04344_),
    .A2(_04345_),
    .A3(_14822_),
    .B1(_04347_),
    .X(_02015_));
 sky130_fd_sc_hd__nand3_1 _20669_ (.A(_04297_),
    .B(_04298_),
    .C(net52),
    .Y(_02016_));
 sky130_vsdinv _20670_ (.A(\count_cycle[27] ),
    .Y(_02019_));
 sky130_fd_sc_hd__and2_1 _20671_ (.A(_04299_),
    .B(_13635_),
    .X(_04348_));
 sky130_fd_sc_hd__a221oi_2 _20672_ (.A1(\count_instr[59] ),
    .A2(_04177_),
    .B1(\count_instr[27] ),
    .B2(_15178_),
    .C1(_04348_),
    .Y(_02020_));
 sky130_fd_sc_hd__and2_1 _20673_ (.A(_14137_),
    .B(\timer[27] ),
    .X(_04349_));
 sky130_fd_sc_hd__a221oi_2 _20674_ (.A1(\irq_mask[27] ),
    .A2(_04264_),
    .B1(\cpuregs_rs1[27] ),
    .B2(_04327_),
    .C1(_04349_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_1 _20675_ (.A(\reg_pc[27] ),
    .B(_14623_),
    .Y(_04350_));
 sky130_fd_sc_hd__and2_1 _20676_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .X(_04351_));
 sky130_fd_sc_hd__nor2_2 _20677_ (.A(_04350_),
    .B(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__and2_1 _20678_ (.A(\reg_pc[26] ),
    .B(_14620_),
    .X(_04353_));
 sky130_fd_sc_hd__or2b_1 _20679_ (.A(_04353_),
    .B_N(_04344_),
    .X(_04354_));
 sky130_fd_sc_hd__o21a_1 _20680_ (.A1(_04352_),
    .A2(_04354_),
    .B1(_14717_),
    .X(_04355_));
 sky130_fd_sc_hd__nand2_1 _20681_ (.A(_04354_),
    .B(_04352_),
    .Y(_04356_));
 sky130_fd_sc_hd__o22ai_1 _20682_ (.A1(_02017_),
    .A2(_04216_),
    .B1(_04217_),
    .B2(_02023_),
    .Y(_04357_));
 sky130_fd_sc_hd__a221o_1 _20683_ (.A1(_14827_),
    .A2(_02018_),
    .B1(_04355_),
    .B2(_04356_),
    .C1(_04357_),
    .X(_02024_));
 sky130_fd_sc_hd__nand3_1 _20684_ (.A(_14818_),
    .B(_15177_),
    .C(net53),
    .Y(_02025_));
 sky130_vsdinv _20685_ (.A(_13691_),
    .Y(_02028_));
 sky130_fd_sc_hd__and2_1 _20686_ (.A(_04299_),
    .B(_13640_),
    .X(_04358_));
 sky130_fd_sc_hd__a221oi_2 _20687_ (.A1(\count_instr[60] ),
    .A2(_04177_),
    .B1(\count_instr[28] ),
    .B2(_15178_),
    .C1(_04358_),
    .Y(_02029_));
 sky130_fd_sc_hd__and2_1 _20688_ (.A(_14137_),
    .B(\timer[28] ),
    .X(_04359_));
 sky130_fd_sc_hd__a221oi_2 _20689_ (.A1(\irq_mask[28] ),
    .A2(_04264_),
    .B1(\cpuregs_rs1[28] ),
    .B2(_04327_),
    .C1(_04359_),
    .Y(_02031_));
 sky130_fd_sc_hd__and2_1 _20690_ (.A(\reg_pc[28] ),
    .B(_14625_),
    .X(_04360_));
 sky130_fd_sc_hd__nand2_1 _20691_ (.A(_04343_),
    .B(_04352_),
    .Y(_04361_));
 sky130_fd_sc_hd__o211a_1 _20692_ (.A1(_13170_),
    .A2(_14623_),
    .B1(\reg_pc[26] ),
    .C1(_14620_),
    .X(_04362_));
 sky130_fd_sc_hd__nor2_1 _20693_ (.A(_04351_),
    .B(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__o21ai_1 _20694_ (.A1(_04361_),
    .A2(_04342_),
    .B1(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__nor2_2 _20695_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .Y(_04365_));
 sky130_vsdinv _20696_ (.A(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand3b_1 _20697_ (.A_N(_04360_),
    .B(_04364_),
    .C(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__o221ai_2 _20698_ (.A1(_04360_),
    .A2(_04365_),
    .B1(_04361_),
    .B2(_04342_),
    .C1(_04363_),
    .Y(_04368_));
 sky130_fd_sc_hd__o2bb2ai_2 _20699_ (.A1_N(_14713_),
    .A2_N(_02027_),
    .B1(_02032_),
    .B2(_04217_),
    .Y(_04369_));
 sky130_fd_sc_hd__and2b_1 _20700_ (.A_N(_02026_),
    .B(_13092_),
    .X(_04370_));
 sky130_fd_sc_hd__a311o_2 _20701_ (.A1(_04367_),
    .A2(_04368_),
    .A3(_14718_),
    .B1(_04369_),
    .C1(_04370_),
    .X(_02033_));
 sky130_fd_sc_hd__nand3_1 _20702_ (.A(_14818_),
    .B(_15177_),
    .C(net54),
    .Y(_02034_));
 sky130_vsdinv _20703_ (.A(\count_cycle[29] ),
    .Y(_02037_));
 sky130_fd_sc_hd__and2_1 _20704_ (.A(\count_instr[61] ),
    .B(_04167_),
    .X(_04371_));
 sky130_fd_sc_hd__a221oi_2 _20705_ (.A1(\count_instr[29] ),
    .A2(_14182_),
    .B1(_04240_),
    .B2(\count_cycle[61] ),
    .C1(_04371_),
    .Y(_02038_));
 sky130_fd_sc_hd__and2_1 _20706_ (.A(\irq_mask[29] ),
    .B(_04252_),
    .X(_04372_));
 sky130_fd_sc_hd__a221oi_2 _20707_ (.A1(_14138_),
    .A2(\timer[29] ),
    .B1(\cpuregs_rs1[29] ),
    .B2(_04327_),
    .C1(_04372_),
    .Y(_02040_));
 sky130_fd_sc_hd__a2bb2oi_4 _20708_ (.A1_N(_02041_),
    .A2_N(_15197_),
    .B1(_13548_),
    .B2(_02036_),
    .Y(_04373_));
 sky130_fd_sc_hd__and2_1 _20709_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .X(_04374_));
 sky130_fd_sc_hd__nor2_2 _20710_ (.A(_13159_),
    .B(\decoded_imm[29] ),
    .Y(_04375_));
 sky130_fd_sc_hd__a21oi_2 _20711_ (.A1(_04364_),
    .A2(_04366_),
    .B1(_04360_),
    .Y(_04376_));
 sky130_fd_sc_hd__nor3_1 _20712_ (.A(_04374_),
    .B(_04375_),
    .C(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__o21ai_1 _20713_ (.A1(_04374_),
    .A2(_04375_),
    .B1(_04376_),
    .Y(_04378_));
 sky130_fd_sc_hd__nand3b_2 _20714_ (.A_N(_04377_),
    .B(_04092_),
    .C(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__o211ai_2 _20715_ (.A1(_15181_),
    .A2(_02035_),
    .B1(_04373_),
    .C1(_04379_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand3_1 _20716_ (.A(_14818_),
    .B(_15177_),
    .C(net497),
    .Y(_02043_));
 sky130_vsdinv _20717_ (.A(\count_cycle[30] ),
    .Y(_02046_));
 sky130_fd_sc_hd__and2_1 _20718_ (.A(\count_instr[30] ),
    .B(instr_rdinstr),
    .X(_04380_));
 sky130_fd_sc_hd__a221oi_2 _20719_ (.A1(\count_instr[62] ),
    .A2(_04177_),
    .B1(_04240_),
    .B2(\count_cycle[62] ),
    .C1(_04380_),
    .Y(_02047_));
 sky130_fd_sc_hd__and2_1 _20720_ (.A(_14137_),
    .B(\timer[30] ),
    .X(_04381_));
 sky130_fd_sc_hd__a221oi_2 _20721_ (.A1(\irq_mask[30] ),
    .A2(_12914_),
    .B1(\cpuregs_rs1[30] ),
    .B2(_04327_),
    .C1(_04381_),
    .Y(_02049_));
 sky130_fd_sc_hd__xor2_1 _20722_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .X(_04382_));
 sky130_fd_sc_hd__o21bai_1 _20723_ (.A1(_04375_),
    .A2(_04376_),
    .B1_N(_04374_),
    .Y(_04383_));
 sky130_fd_sc_hd__o21a_1 _20724_ (.A1(_04382_),
    .A2(_04383_),
    .B1(_14717_),
    .X(_04384_));
 sky130_fd_sc_hd__nand2_1 _20725_ (.A(_04383_),
    .B(_04382_),
    .Y(_04385_));
 sky130_fd_sc_hd__and2b_1 _20726_ (.A_N(_02044_),
    .B(_12652_),
    .X(_04386_));
 sky130_fd_sc_hd__o2bb2ai_2 _20727_ (.A1_N(_15167_),
    .A2_N(_02045_),
    .B1(_02050_),
    .B2(_15197_),
    .Y(_04387_));
 sky130_fd_sc_hd__a211o_1 _20728_ (.A1(_04384_),
    .A2(_04385_),
    .B1(_04386_),
    .C1(_04387_),
    .X(_02051_));
 sky130_fd_sc_hd__nand3_1 _20729_ (.A(_14818_),
    .B(_15177_),
    .C(net57),
    .Y(_02052_));
 sky130_vsdinv _20730_ (.A(_13594_),
    .Y(_02055_));
 sky130_fd_sc_hd__and2_1 _20731_ (.A(\count_instr[63] ),
    .B(_04167_),
    .X(_04388_));
 sky130_fd_sc_hd__a221oi_2 _20732_ (.A1(\count_instr[31] ),
    .A2(_14182_),
    .B1(_14185_),
    .B2(\count_cycle[63] ),
    .C1(_04388_),
    .Y(_02056_));
 sky130_fd_sc_hd__and2_1 _20733_ (.A(\irq_mask[31] ),
    .B(_12908_),
    .X(_04389_));
 sky130_fd_sc_hd__a221oi_2 _20734_ (.A1(_14138_),
    .A2(\timer[31] ),
    .B1(\cpuregs_rs1[31] ),
    .B2(_15190_),
    .C1(_04389_),
    .Y(_02058_));
 sky130_fd_sc_hd__and2_1 _20735_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .X(_04390_));
 sky130_vsdinv _20736_ (.A(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__xnor2_1 _20737_ (.A(\reg_pc[31] ),
    .B(\decoded_imm[31] ),
    .Y(_04392_));
 sky130_fd_sc_hd__a21oi_1 _20738_ (.A1(_04385_),
    .A2(_04391_),
    .B1(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__a31o_1 _20739_ (.A1(_04385_),
    .A2(_04391_),
    .A3(_04392_),
    .B1(_12812_),
    .X(_04394_));
 sky130_fd_sc_hd__nand2_1 _20740_ (.A(_04125_),
    .B(_02054_),
    .Y(_04395_));
 sky130_fd_sc_hd__o221ai_2 _20741_ (.A1(_02053_),
    .A2(_04216_),
    .B1(_02059_),
    .B2(_04217_),
    .C1(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__o21bai_2 _20742_ (.A1(_04393_),
    .A2(_04394_),
    .B1_N(_04396_),
    .Y(_02060_));
 sky130_fd_sc_hd__nand3b_1 _20743_ (.A_N(\decoded_rd[4] ),
    .B(_12771_),
    .C(_12873_),
    .Y(_02061_));
 sky130_vsdinv _20744_ (.A(instr_jalr),
    .Y(_02063_));
 sky130_fd_sc_hd__o21bai_1 _20745_ (.A1(_02064_),
    .A2(_12813_),
    .B1_N(_12917_),
    .Y(_02065_));
 sky130_fd_sc_hd__o211a_1 _20746_ (.A1(_13558_),
    .A2(_13564_),
    .B1(_00309_),
    .C1(_12774_),
    .X(_02066_));
 sky130_fd_sc_hd__and3_1 _20747_ (.A(_12850_),
    .B(_15182_),
    .C(_12660_),
    .X(_02067_));
 sky130_fd_sc_hd__and2_1 _20748_ (.A(_12979_),
    .B(_00343_),
    .X(_04397_));
 sky130_fd_sc_hd__o211ai_2 _20749_ (.A1(_12813_),
    .A2(_04397_),
    .B1(_15184_),
    .C1(_15181_),
    .Y(_02068_));
 sky130_fd_sc_hd__o21a_2 _20750_ (.A1(_14536_),
    .A2(_13736_),
    .B1(_12873_),
    .X(_02069_));
 sky130_vsdinv _20751_ (.A(_12863_),
    .Y(_04398_));
 sky130_fd_sc_hd__buf_6 _20752_ (.A(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__buf_6 _20753_ (.A(_13455_),
    .X(_04400_));
 sky130_fd_sc_hd__nand3b_2 _20754_ (.A_N(_12663_),
    .B(_12858_),
    .C(_02070_),
    .Y(_04401_));
 sky130_fd_sc_hd__o221ai_1 _20755_ (.A1(_04399_),
    .A2(_14535_),
    .B1(_04400_),
    .B2(_12755_),
    .C1(_04401_),
    .Y(_02071_));
 sky130_fd_sc_hd__clkbuf_4 _20756_ (.A(_13455_),
    .X(_04402_));
 sky130_fd_sc_hd__buf_2 _20757_ (.A(_13735_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_4 _20758_ (.A(_12857_),
    .X(_04404_));
 sky130_fd_sc_hd__a32oi_1 _20759_ (.A1(_04403_),
    .A2(_04404_),
    .A3(_01465_),
    .B1(_12864_),
    .B2(\reg_next_pc[1] ),
    .Y(_04405_));
 sky130_fd_sc_hd__o21ai_1 _20760_ (.A1(_04402_),
    .A2(_12757_),
    .B1(_04405_),
    .Y(_02072_));
 sky130_vsdinv _20761_ (.A(_13249_),
    .Y(_02073_));
 sky130_fd_sc_hd__and2b_1 _20762_ (.A_N(latched_branch),
    .B(latched_store),
    .X(_04406_));
 sky130_fd_sc_hd__buf_2 _20763_ (.A(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__nand3b_2 _20764_ (.A_N(\irq_mask[2] ),
    .B(_12862_),
    .C(\irq_pending[2] ),
    .Y(_04408_));
 sky130_vsdinv _20765_ (.A(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__a221o_1 _20766_ (.A1(_15011_),
    .A2(\reg_next_pc[2] ),
    .B1(_00293_),
    .B2(_04407_),
    .C1(_04409_),
    .X(_02074_));
 sky130_fd_sc_hd__xor2_1 _20767_ (.A(_13246_),
    .B(_13249_),
    .X(_02075_));
 sky130_fd_sc_hd__nand3b_1 _20768_ (.A_N(\irq_mask[3] ),
    .B(_12862_),
    .C(\irq_pending[3] ),
    .Y(_04410_));
 sky130_vsdinv _20769_ (.A(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__a221o_1 _20770_ (.A1(_15011_),
    .A2(\reg_next_pc[3] ),
    .B1(_01468_),
    .B2(_04407_),
    .C1(_04411_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_1 _20771_ (.A(_13246_),
    .B(_13249_),
    .Y(_04412_));
 sky130_fd_sc_hd__xnor2_1 _20772_ (.A(_13244_),
    .B(_04412_),
    .Y(_02077_));
 sky130_fd_sc_hd__clkbuf_2 _20773_ (.A(latched_branch),
    .X(_04413_));
 sky130_fd_sc_hd__nand3b_2 _20774_ (.A_N(_04413_),
    .B(_12858_),
    .C(_01472_),
    .Y(_04414_));
 sky130_fd_sc_hd__o221ai_4 _20775_ (.A1(_04399_),
    .A2(_01471_),
    .B1(_04400_),
    .B2(_12737_),
    .C1(_04414_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand3_2 _20776_ (.A(_13244_),
    .B(_13246_),
    .C(_13249_),
    .Y(_04415_));
 sky130_fd_sc_hd__xnor2_1 _20777_ (.A(_13241_),
    .B(_04415_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand3b_2 _20778_ (.A_N(_04413_),
    .B(_12858_),
    .C(_01476_),
    .Y(_04416_));
 sky130_fd_sc_hd__o221ai_4 _20779_ (.A1(_04399_),
    .A2(_13147_),
    .B1(_04400_),
    .B2(_12741_),
    .C1(_04416_),
    .Y(_02080_));
 sky130_fd_sc_hd__and4_2 _20780_ (.A(_13241_),
    .B(_13244_),
    .C(_13246_),
    .D(\reg_pc[2] ),
    .X(_04417_));
 sky130_fd_sc_hd__xor2_1 _20781_ (.A(_13237_),
    .B(_04417_),
    .X(_02081_));
 sky130_fd_sc_hd__nand3b_1 _20782_ (.A_N(\irq_mask[6] ),
    .B(_12862_),
    .C(\irq_pending[6] ),
    .Y(_04418_));
 sky130_vsdinv _20783_ (.A(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__a221o_1 _20784_ (.A1(_15011_),
    .A2(\reg_next_pc[6] ),
    .B1(_01479_),
    .B2(_04407_),
    .C1(_04419_),
    .X(_02082_));
 sky130_fd_sc_hd__nand3b_2 _20785_ (.A_N(_04415_),
    .B(_13237_),
    .C(_13241_),
    .Y(_04420_));
 sky130_fd_sc_hd__xnor2_1 _20786_ (.A(\reg_pc[7] ),
    .B(_04420_),
    .Y(_02083_));
 sky130_fd_sc_hd__a32oi_2 _20787_ (.A1(_04403_),
    .A2(_04404_),
    .A3(_01482_),
    .B1(_12864_),
    .B2(\reg_next_pc[7] ),
    .Y(_04421_));
 sky130_fd_sc_hd__o21ai_2 _20788_ (.A1(_04402_),
    .A2(_12739_),
    .B1(_04421_),
    .Y(_02084_));
 sky130_fd_sc_hd__nand3_4 _20789_ (.A(_04417_),
    .B(\reg_pc[7] ),
    .C(_13237_),
    .Y(_04422_));
 sky130_fd_sc_hd__xor2_1 _20790_ (.A(_13233_),
    .B(_04422_),
    .X(_02085_));
 sky130_fd_sc_hd__clkbuf_2 _20791_ (.A(_12861_),
    .X(_04423_));
 sky130_fd_sc_hd__nand3b_1 _20792_ (.A_N(\irq_mask[8] ),
    .B(_04423_),
    .C(\irq_pending[8] ),
    .Y(_04424_));
 sky130_vsdinv _20793_ (.A(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__a221o_1 _20794_ (.A1(_15011_),
    .A2(\reg_next_pc[8] ),
    .B1(_01485_),
    .B2(_04407_),
    .C1(_04425_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_2 _20795_ (.A(_13233_),
    .B(_04422_),
    .Y(_04426_));
 sky130_fd_sc_hd__xor2_1 _20796_ (.A(_13229_),
    .B(_04426_),
    .X(_02087_));
 sky130_fd_sc_hd__a32oi_2 _20797_ (.A1(_04403_),
    .A2(_04404_),
    .A3(_01488_),
    .B1(_12864_),
    .B2(\reg_next_pc[9] ),
    .Y(_04427_));
 sky130_fd_sc_hd__o21ai_2 _20798_ (.A1(_04402_),
    .A2(_12723_),
    .B1(_04427_),
    .Y(_02088_));
 sky130_fd_sc_hd__nor3b_4 _20799_ (.A(_13233_),
    .B(_04422_),
    .C_N(_13229_),
    .Y(_04428_));
 sky130_fd_sc_hd__xor2_1 _20800_ (.A(_13226_),
    .B(_04428_),
    .X(_02089_));
 sky130_fd_sc_hd__nand3b_1 _20801_ (.A_N(\irq_mask[10] ),
    .B(_04423_),
    .C(\irq_pending[10] ),
    .Y(_04429_));
 sky130_vsdinv _20802_ (.A(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__a221o_1 _20803_ (.A1(_15011_),
    .A2(\reg_next_pc[10] ),
    .B1(_01491_),
    .B2(_04407_),
    .C1(_04430_),
    .X(_02090_));
 sky130_fd_sc_hd__nand3_1 _20804_ (.A(_04426_),
    .B(_13226_),
    .C(_13229_),
    .Y(_04431_));
 sky130_fd_sc_hd__xnor2_1 _20805_ (.A(_13223_),
    .B(_04431_),
    .Y(_02091_));
 sky130_fd_sc_hd__a32oi_2 _20806_ (.A1(_04403_),
    .A2(_12857_),
    .A3(_01494_),
    .B1(_12864_),
    .B2(\reg_next_pc[11] ),
    .Y(_04432_));
 sky130_fd_sc_hd__o21ai_2 _20807_ (.A1(_04402_),
    .A2(_12721_),
    .B1(_04432_),
    .Y(_02092_));
 sky130_fd_sc_hd__nand3_4 _20808_ (.A(_04428_),
    .B(_13223_),
    .C(_13226_),
    .Y(_04433_));
 sky130_fd_sc_hd__xor2_1 _20809_ (.A(_13220_),
    .B(_04433_),
    .X(_02093_));
 sky130_fd_sc_hd__buf_2 _20810_ (.A(_12863_),
    .X(_04434_));
 sky130_fd_sc_hd__buf_2 _20811_ (.A(_04406_),
    .X(_04435_));
 sky130_fd_sc_hd__nand3b_1 _20812_ (.A_N(\irq_mask[12] ),
    .B(_04423_),
    .C(\irq_pending[12] ),
    .Y(_04436_));
 sky130_vsdinv _20813_ (.A(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__a221o_1 _20814_ (.A1(_04434_),
    .A2(\reg_next_pc[12] ),
    .B1(_01497_),
    .B2(_04435_),
    .C1(_04437_),
    .X(_02094_));
 sky130_fd_sc_hd__nor2_4 _20815_ (.A(_13220_),
    .B(_04433_),
    .Y(_04438_));
 sky130_fd_sc_hd__xor2_1 _20816_ (.A(_13215_),
    .B(_04438_),
    .X(_02095_));
 sky130_fd_sc_hd__buf_2 _20817_ (.A(_12857_),
    .X(_04439_));
 sky130_fd_sc_hd__nand3b_2 _20818_ (.A_N(_04413_),
    .B(_04439_),
    .C(_01500_),
    .Y(_04440_));
 sky130_fd_sc_hd__o221ai_4 _20819_ (.A1(_04399_),
    .A2(_13134_),
    .B1(_04400_),
    .B2(_12714_),
    .C1(_04440_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor3b_4 _20820_ (.A(_13220_),
    .B(_04433_),
    .C_N(_13215_),
    .Y(_04441_));
 sky130_fd_sc_hd__xor2_1 _20821_ (.A(_13213_),
    .B(_04441_),
    .X(_02097_));
 sky130_fd_sc_hd__nand3b_4 _20822_ (.A_N(\irq_mask[14] ),
    .B(_12862_),
    .C(\irq_pending[14] ),
    .Y(_04442_));
 sky130_fd_sc_hd__nand3b_2 _20823_ (.A_N(_12663_),
    .B(_12858_),
    .C(_01503_),
    .Y(_04443_));
 sky130_fd_sc_hd__o211ai_4 _20824_ (.A1(_04399_),
    .A2(_13132_),
    .B1(_04442_),
    .C1(_04443_),
    .Y(_02098_));
 sky130_fd_sc_hd__nand3_1 _20825_ (.A(_04438_),
    .B(_13213_),
    .C(_13215_),
    .Y(_04444_));
 sky130_fd_sc_hd__xnor2_1 _20826_ (.A(_13208_),
    .B(_04444_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand3b_2 _20827_ (.A_N(_04413_),
    .B(_04439_),
    .C(_01506_),
    .Y(_04445_));
 sky130_fd_sc_hd__o221ai_4 _20828_ (.A1(_04399_),
    .A2(_13130_),
    .B1(_04400_),
    .B2(_12712_),
    .C1(_04445_),
    .Y(_02100_));
 sky130_vsdinv _20829_ (.A(_13205_),
    .Y(_04446_));
 sky130_fd_sc_hd__nand3_2 _20830_ (.A(_04441_),
    .B(_13208_),
    .C(_13213_),
    .Y(_04447_));
 sky130_fd_sc_hd__xor2_1 _20831_ (.A(_04446_),
    .B(_04447_),
    .X(_02101_));
 sky130_fd_sc_hd__nand3b_1 _20832_ (.A_N(\irq_mask[16] ),
    .B(_04423_),
    .C(\irq_pending[16] ),
    .Y(_04448_));
 sky130_vsdinv _20833_ (.A(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__a221o_1 _20834_ (.A1(_04434_),
    .A2(\reg_next_pc[16] ),
    .B1(_01509_),
    .B2(_04435_),
    .C1(_04449_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_2 _20835_ (.A(_04446_),
    .B(_04447_),
    .Y(_04450_));
 sky130_fd_sc_hd__xor2_1 _20836_ (.A(_13203_),
    .B(_04450_),
    .X(_02103_));
 sky130_fd_sc_hd__buf_4 _20837_ (.A(_04398_),
    .X(_04451_));
 sky130_fd_sc_hd__nand3b_2 _20838_ (.A_N(_04413_),
    .B(_04439_),
    .C(_01512_),
    .Y(_04452_));
 sky130_fd_sc_hd__o221ai_4 _20839_ (.A1(_04451_),
    .A2(_13125_),
    .B1(_04400_),
    .B2(_12766_),
    .C1(_04452_),
    .Y(_02104_));
 sky130_fd_sc_hd__and4_1 _20840_ (.A(_04426_),
    .B(_13223_),
    .C(_13226_),
    .D(_13229_),
    .X(_04453_));
 sky130_fd_sc_hd__and4_1 _20841_ (.A(_04453_),
    .B(_13213_),
    .C(_13215_),
    .D(\reg_pc[12] ),
    .X(_04454_));
 sky130_fd_sc_hd__and4_2 _20842_ (.A(_04454_),
    .B(_13203_),
    .C(_13205_),
    .D(_13208_),
    .X(_04455_));
 sky130_fd_sc_hd__xor2_1 _20843_ (.A(_13199_),
    .B(_04455_),
    .X(_02105_));
 sky130_fd_sc_hd__nand3b_1 _20844_ (.A_N(\irq_mask[18] ),
    .B(_04423_),
    .C(\irq_pending[18] ),
    .Y(_04456_));
 sky130_vsdinv _20845_ (.A(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__a221o_1 _20846_ (.A1(_04434_),
    .A2(\reg_next_pc[18] ),
    .B1(_01515_),
    .B2(_04435_),
    .C1(_04457_),
    .X(_02106_));
 sky130_fd_sc_hd__nand3_1 _20847_ (.A(_04450_),
    .B(_13199_),
    .C(_13203_),
    .Y(_04458_));
 sky130_fd_sc_hd__xnor2_1 _20848_ (.A(_13194_),
    .B(_04458_),
    .Y(_02107_));
 sky130_fd_sc_hd__clkbuf_4 _20849_ (.A(_13455_),
    .X(_04459_));
 sky130_fd_sc_hd__nand3b_2 _20850_ (.A_N(_04413_),
    .B(_04439_),
    .C(_01518_),
    .Y(_04460_));
 sky130_fd_sc_hd__o221ai_4 _20851_ (.A1(_04451_),
    .A2(_13122_),
    .B1(_04459_),
    .B2(_12764_),
    .C1(_04460_),
    .Y(_02108_));
 sky130_fd_sc_hd__and4_2 _20852_ (.A(_04450_),
    .B(_13194_),
    .C(_13199_),
    .D(_13203_),
    .X(_04461_));
 sky130_fd_sc_hd__xor2_1 _20853_ (.A(_13192_),
    .B(_04461_),
    .X(_02109_));
 sky130_fd_sc_hd__nand3b_1 _20854_ (.A_N(_14537_),
    .B(_04439_),
    .C(_01521_),
    .Y(_04462_));
 sky130_fd_sc_hd__o221ai_1 _20855_ (.A1(_04451_),
    .A2(_13120_),
    .B1(_04459_),
    .B2(_12731_),
    .C1(_04462_),
    .Y(_02110_));
 sky130_fd_sc_hd__and4_1 _20856_ (.A(_04455_),
    .B(_13192_),
    .C(_13194_),
    .D(\reg_pc[18] ),
    .X(_04463_));
 sky130_fd_sc_hd__xor2_1 _20857_ (.A(_13189_),
    .B(_04463_),
    .X(_02111_));
 sky130_fd_sc_hd__nand3b_1 _20858_ (.A_N(_14537_),
    .B(_04439_),
    .C(_01524_),
    .Y(_04464_));
 sky130_fd_sc_hd__o221ai_1 _20859_ (.A1(_04451_),
    .A2(_13117_),
    .B1(_04459_),
    .B2(_12727_),
    .C1(_04464_),
    .Y(_02112_));
 sky130_fd_sc_hd__and4_1 _20860_ (.A(_04438_),
    .B(_13208_),
    .C(\reg_pc[14] ),
    .D(\reg_pc[13] ),
    .X(_04465_));
 sky130_fd_sc_hd__and4_1 _20861_ (.A(_04465_),
    .B(\reg_pc[18] ),
    .C(\reg_pc[17] ),
    .D(_13205_),
    .X(_04466_));
 sky130_fd_sc_hd__and4_2 _20862_ (.A(_04466_),
    .B(_13189_),
    .C(_13192_),
    .D(_13194_),
    .X(_04467_));
 sky130_fd_sc_hd__xor2_1 _20863_ (.A(_13186_),
    .B(_04467_),
    .X(_02113_));
 sky130_fd_sc_hd__nand3b_1 _20864_ (.A_N(\irq_mask[22] ),
    .B(_04423_),
    .C(\irq_pending[22] ),
    .Y(_04468_));
 sky130_vsdinv _20865_ (.A(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__a221o_1 _20866_ (.A1(_04434_),
    .A2(\reg_next_pc[22] ),
    .B1(_01527_),
    .B2(_04435_),
    .C1(_04469_),
    .X(_02114_));
 sky130_fd_sc_hd__and4_1 _20867_ (.A(_04461_),
    .B(_13186_),
    .C(_13189_),
    .D(_13192_),
    .X(_04470_));
 sky130_fd_sc_hd__xor2_1 _20868_ (.A(_13182_),
    .B(_04470_),
    .X(_02115_));
 sky130_fd_sc_hd__nand3b_1 _20869_ (.A_N(\irq_mask[23] ),
    .B(_12861_),
    .C(\irq_pending[23] ),
    .Y(_04471_));
 sky130_vsdinv _20870_ (.A(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__a221o_1 _20871_ (.A1(_04434_),
    .A2(\reg_next_pc[23] ),
    .B1(_01530_),
    .B2(_04435_),
    .C1(_04472_),
    .X(_02116_));
 sky130_vsdinv _20872_ (.A(\reg_pc[24] ),
    .Y(_04473_));
 sky130_fd_sc_hd__nand3_4 _20873_ (.A(_04467_),
    .B(_13182_),
    .C(_13186_),
    .Y(_04474_));
 sky130_fd_sc_hd__xor2_1 _20874_ (.A(_04473_),
    .B(_04474_),
    .X(_02117_));
 sky130_fd_sc_hd__nand3b_2 _20875_ (.A_N(_14537_),
    .B(_04404_),
    .C(_01533_),
    .Y(_04475_));
 sky130_fd_sc_hd__o221ai_2 _20876_ (.A1(_04451_),
    .A2(_13110_),
    .B1(_04459_),
    .B2(_12749_),
    .C1(_04475_),
    .Y(_02118_));
 sky130_fd_sc_hd__nor2_2 _20877_ (.A(_04473_),
    .B(_04474_),
    .Y(_04476_));
 sky130_fd_sc_hd__xor2_1 _20878_ (.A(_13175_),
    .B(_04476_),
    .X(_02119_));
 sky130_fd_sc_hd__nand3b_1 _20879_ (.A_N(\irq_mask[25] ),
    .B(_12861_),
    .C(\irq_pending[25] ),
    .Y(_04477_));
 sky130_vsdinv _20880_ (.A(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__a221o_1 _20881_ (.A1(_04434_),
    .A2(\reg_next_pc[25] ),
    .B1(_01536_),
    .B2(_04435_),
    .C1(_04478_),
    .X(_02120_));
 sky130_fd_sc_hd__nor3b_4 _20882_ (.A(_04473_),
    .B(_04474_),
    .C_N(_13175_),
    .Y(_04479_));
 sky130_fd_sc_hd__xor2_1 _20883_ (.A(_13173_),
    .B(_04479_),
    .X(_02121_));
 sky130_fd_sc_hd__nand3b_2 _20884_ (.A_N(_14537_),
    .B(_04404_),
    .C(_01539_),
    .Y(_04480_));
 sky130_fd_sc_hd__o221ai_2 _20885_ (.A1(_04451_),
    .A2(_13107_),
    .B1(_04459_),
    .B2(_12747_),
    .C1(_04480_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand3_1 _20886_ (.A(_04476_),
    .B(_13173_),
    .C(_13175_),
    .Y(_04481_));
 sky130_fd_sc_hd__xnor2_1 _20887_ (.A(_13170_),
    .B(_04481_),
    .Y(_02123_));
 sky130_fd_sc_hd__a32oi_1 _20888_ (.A1(_04403_),
    .A2(_12857_),
    .A3(_01542_),
    .B1(_12878_),
    .B2(\reg_next_pc[27] ),
    .Y(_04482_));
 sky130_fd_sc_hd__o31ai_1 _20889_ (.A1(_04402_),
    .A2(\irq_mask[27] ),
    .A3(_12743_),
    .B1(_04482_),
    .Y(_02124_));
 sky130_vsdinv _20890_ (.A(\reg_pc[28] ),
    .Y(_04483_));
 sky130_fd_sc_hd__nand3_2 _20891_ (.A(_04479_),
    .B(_13170_),
    .C(_13173_),
    .Y(_04484_));
 sky130_fd_sc_hd__xor2_1 _20892_ (.A(_04483_),
    .B(_04484_),
    .X(_02125_));
 sky130_fd_sc_hd__nand3b_1 _20893_ (.A_N(_14537_),
    .B(_04404_),
    .C(_01545_),
    .Y(_04485_));
 sky130_fd_sc_hd__o221ai_1 _20894_ (.A1(_04398_),
    .A2(_13104_),
    .B1(_04459_),
    .B2(_12706_),
    .C1(_04485_),
    .Y(_02126_));
 sky130_fd_sc_hd__nor2_2 _20895_ (.A(_04483_),
    .B(_04484_),
    .Y(_04486_));
 sky130_fd_sc_hd__xor2_1 _20896_ (.A(_13159_),
    .B(_04486_),
    .X(_02127_));
 sky130_fd_sc_hd__a32oi_1 _20897_ (.A1(_04403_),
    .A2(_12857_),
    .A3(_01548_),
    .B1(_12878_),
    .B2(\reg_next_pc[29] ),
    .Y(_04487_));
 sky130_fd_sc_hd__o21ai_1 _20898_ (.A1(_04402_),
    .A2(_12702_),
    .B1(_04487_),
    .Y(_02128_));
 sky130_fd_sc_hd__and4_1 _20899_ (.A(_04463_),
    .B(_13182_),
    .C(_13186_),
    .D(_13189_),
    .X(_04488_));
 sky130_fd_sc_hd__and4_1 _20900_ (.A(_04488_),
    .B(_13173_),
    .C(_13175_),
    .D(\reg_pc[24] ),
    .X(_04489_));
 sky130_fd_sc_hd__and4_1 _20901_ (.A(_04489_),
    .B(_13159_),
    .C(\reg_pc[28] ),
    .D(_13170_),
    .X(_04490_));
 sky130_fd_sc_hd__xor2_1 _20902_ (.A(\reg_pc[30] ),
    .B(_04490_),
    .X(_02129_));
 sky130_fd_sc_hd__o2bb2ai_1 _20903_ (.A1_N(_12878_),
    .A2_N(\reg_next_pc[30] ),
    .B1(_13455_),
    .B2(_12704_),
    .Y(_04491_));
 sky130_fd_sc_hd__a21o_1 _20904_ (.A1(_01551_),
    .A2(_04407_),
    .B1(_04491_),
    .X(_02130_));
 sky130_fd_sc_hd__nand3_1 _20905_ (.A(_04486_),
    .B(\reg_pc[30] ),
    .C(_13159_),
    .Y(_04492_));
 sky130_fd_sc_hd__xor2_1 _20906_ (.A(_13155_),
    .B(_04492_),
    .X(_02131_));
 sky130_fd_sc_hd__nand3b_1 _20907_ (.A_N(\irq_mask[31] ),
    .B(_12861_),
    .C(\irq_pending[31] ),
    .Y(_04493_));
 sky130_vsdinv _20908_ (.A(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__a221o_1 _20909_ (.A1(_12864_),
    .A2(\reg_next_pc[31] ),
    .B1(_01554_),
    .B2(_04406_),
    .C1(_04494_),
    .X(_02132_));
 sky130_fd_sc_hd__or2_2 _20910_ (.A(instr_xor),
    .B(instr_xori),
    .X(_04495_));
 sky130_fd_sc_hd__buf_2 _20911_ (.A(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__nor3b_2 _20912_ (.A(is_compare),
    .B(_04496_),
    .C_N(_12828_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor2_4 _20913_ (.A(instr_sll),
    .B(instr_slli),
    .Y(_04498_));
 sky130_fd_sc_hd__nor2_4 _20914_ (.A(instr_or),
    .B(instr_ori),
    .Y(_04499_));
 sky130_fd_sc_hd__clkbuf_2 _20915_ (.A(_04499_),
    .X(_04500_));
 sky130_fd_sc_hd__clkbuf_4 _20916_ (.A(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__nor2_4 _20917_ (.A(instr_and),
    .B(instr_andi),
    .Y(_04502_));
 sky130_fd_sc_hd__clkbuf_2 _20918_ (.A(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__and4_4 _20919_ (.A(_04497_),
    .B(_04498_),
    .C(_04501_),
    .D(_04503_),
    .X(_02133_));
 sky130_fd_sc_hd__o21ai_1 _20920_ (.A1(_15170_),
    .A2(_04503_),
    .B1(_04501_),
    .Y(_04504_));
 sky130_vsdinv _20921_ (.A(_12828_),
    .Y(_04505_));
 sky130_fd_sc_hd__clkbuf_2 _20922_ (.A(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__buf_2 _20923_ (.A(_04506_),
    .X(_04507_));
 sky130_vsdinv _20924_ (.A(_04498_),
    .Y(_04508_));
 sky130_vsdinv _20925_ (.A(_04499_),
    .Y(_04509_));
 sky130_fd_sc_hd__and2b_1 _20926_ (.A_N(_00343_),
    .B(is_compare),
    .X(_04510_));
 sky130_fd_sc_hd__a221o_1 _20927_ (.A1(_04508_),
    .A2(\alu_shl[0] ),
    .B1(_04509_),
    .B2(_14267_),
    .C1(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__a221o_1 _20928_ (.A1(\alu_shr[0] ),
    .A2(_04507_),
    .B1(_02591_),
    .B2(_04496_),
    .C1(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__a21o_1 _20929_ (.A1(_13840_),
    .A2(_04504_),
    .B1(_04512_),
    .X(_02134_));
 sky130_fd_sc_hd__o211ai_1 _20930_ (.A1(_13007_),
    .A2(_13050_),
    .B1(_13837_),
    .C1(_15172_),
    .Y(_04513_));
 sky130_fd_sc_hd__buf_2 _20931_ (.A(_04508_),
    .X(_04514_));
 sky130_fd_sc_hd__clkbuf_4 _20932_ (.A(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__clkbuf_4 _20933_ (.A(_04506_),
    .X(_04516_));
 sky130_fd_sc_hd__buf_2 _20934_ (.A(_04495_),
    .X(_04517_));
 sky130_fd_sc_hd__nor3b_4 _20935_ (.A(_14774_),
    .B(_14775_),
    .C_N(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__a221oi_2 _20936_ (.A1(\alu_shl[1] ),
    .A2(_04515_),
    .B1(_04516_),
    .B2(\alu_shr[1] ),
    .C1(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__o211ai_1 _20937_ (.A1(_14774_),
    .A2(_04501_),
    .B1(_04513_),
    .C1(_04519_),
    .Y(_02135_));
 sky130_fd_sc_hd__clkbuf_2 _20938_ (.A(_04514_),
    .X(_04520_));
 sky130_fd_sc_hd__clkbuf_2 _20939_ (.A(_04496_),
    .X(_04521_));
 sky130_fd_sc_hd__a211oi_2 _20940_ (.A1(_13835_),
    .A2(_14262_),
    .B1(_13012_),
    .C1(_13053_),
    .Y(_04522_));
 sky130_fd_sc_hd__o2bb2ai_1 _20941_ (.A1_N(_04500_),
    .A2_N(_04503_),
    .B1(_13835_),
    .B2(_14262_),
    .Y(_04523_));
 sky130_fd_sc_hd__o2bb2ai_1 _20942_ (.A1_N(\alu_shr[2] ),
    .A2_N(_04516_),
    .B1(_04522_),
    .B2(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__a221o_1 _20943_ (.A1(\alu_shl[2] ),
    .A2(_04520_),
    .B1(_14787_),
    .B2(_04521_),
    .C1(_04524_),
    .X(_02136_));
 sky130_fd_sc_hd__clkbuf_2 _20944_ (.A(_04506_),
    .X(_04525_));
 sky130_fd_sc_hd__a211oi_4 _20945_ (.A1(_13833_),
    .A2(_14260_),
    .B1(_13012_),
    .C1(_13053_),
    .Y(_04526_));
 sky130_fd_sc_hd__o2bb2ai_1 _20946_ (.A1_N(_04500_),
    .A2_N(_04503_),
    .B1(_13833_),
    .B2(_14260_),
    .Y(_04527_));
 sky130_fd_sc_hd__o2bb2ai_1 _20947_ (.A1_N(\alu_shr[3] ),
    .A2_N(_04525_),
    .B1(_04526_),
    .B2(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__a221o_1 _20948_ (.A1(\alu_shl[3] ),
    .A2(_04520_),
    .B1(_14781_),
    .B2(_04521_),
    .C1(_04528_),
    .X(_02137_));
 sky130_fd_sc_hd__buf_2 _20949_ (.A(instr_or),
    .X(_04529_));
 sky130_fd_sc_hd__buf_2 _20950_ (.A(instr_ori),
    .X(_04530_));
 sky130_fd_sc_hd__o22a_1 _20951_ (.A1(_04529_),
    .A2(_04530_),
    .B1(_13831_),
    .B2(_14259_),
    .X(_04531_));
 sky130_fd_sc_hd__o211a_1 _20952_ (.A1(_13007_),
    .A2(_13050_),
    .B1(_13831_),
    .C1(_14259_),
    .X(_04532_));
 sky130_fd_sc_hd__a211o_1 _20953_ (.A1(_04507_),
    .A2(\alu_shr[4] ),
    .B1(_04531_),
    .C1(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__a221o_1 _20954_ (.A1(\alu_shl[4] ),
    .A2(_04520_),
    .B1(_14791_),
    .B2(_04521_),
    .C1(_04533_),
    .X(_02138_));
 sky130_fd_sc_hd__nor2_1 _20955_ (.A(_14776_),
    .B(_14777_),
    .Y(_04534_));
 sky130_fd_sc_hd__a211oi_4 _20956_ (.A1(_13829_),
    .A2(_14257_),
    .B1(_13012_),
    .C1(_13053_),
    .Y(_04535_));
 sky130_fd_sc_hd__o2bb2ai_1 _20957_ (.A1_N(_04500_),
    .A2_N(_04503_),
    .B1(_13829_),
    .B2(_14257_),
    .Y(_04536_));
 sky130_fd_sc_hd__o2bb2ai_1 _20958_ (.A1_N(\alu_shr[5] ),
    .A2_N(_04525_),
    .B1(_04535_),
    .B2(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__a221o_1 _20959_ (.A1(\alu_shl[5] ),
    .A2(_04520_),
    .B1(_04534_),
    .B2(_04521_),
    .C1(_04537_),
    .X(_02139_));
 sky130_vsdinv _20960_ (.A(_14788_),
    .Y(_04538_));
 sky130_fd_sc_hd__buf_2 _20961_ (.A(_04509_),
    .X(_04539_));
 sky130_fd_sc_hd__clkbuf_2 _20962_ (.A(_04505_),
    .X(_04540_));
 sky130_fd_sc_hd__clkbuf_2 _20963_ (.A(instr_and),
    .X(_04541_));
 sky130_fd_sc_hd__clkbuf_2 _20964_ (.A(instr_andi),
    .X(_04542_));
 sky130_fd_sc_hd__o211a_1 _20965_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_13827_),
    .C1(_14256_),
    .X(_04543_));
 sky130_fd_sc_hd__a221o_1 _20966_ (.A1(_04538_),
    .A2(_04539_),
    .B1(_04540_),
    .B2(\alu_shr[6] ),
    .C1(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__a221o_1 _20967_ (.A1(\alu_shl[6] ),
    .A2(_04520_),
    .B1(_14790_),
    .B2(_04521_),
    .C1(_04544_),
    .X(_02140_));
 sky130_fd_sc_hd__clkbuf_2 _20968_ (.A(_04514_),
    .X(_04545_));
 sky130_fd_sc_hd__a211oi_2 _20969_ (.A1(_13825_),
    .A2(_14253_),
    .B1(_13012_),
    .C1(_13053_),
    .Y(_04546_));
 sky130_fd_sc_hd__clkbuf_2 _20970_ (.A(_04502_),
    .X(_04547_));
 sky130_fd_sc_hd__o2bb2ai_1 _20971_ (.A1_N(_04500_),
    .A2_N(_04547_),
    .B1(_13825_),
    .B2(_14253_),
    .Y(_04548_));
 sky130_fd_sc_hd__o2bb2ai_1 _20972_ (.A1_N(\alu_shr[7] ),
    .A2_N(_04525_),
    .B1(_04546_),
    .B2(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__a221o_1 _20973_ (.A1(\alu_shl[7] ),
    .A2(_04545_),
    .B1(_14786_),
    .B2(_04521_),
    .C1(_04549_),
    .X(_02141_));
 sky130_fd_sc_hd__clkbuf_2 _20974_ (.A(_04517_),
    .X(_04550_));
 sky130_fd_sc_hd__o22a_1 _20975_ (.A1(_04529_),
    .A2(_04530_),
    .B1(_13823_),
    .B2(_14251_),
    .X(_04551_));
 sky130_fd_sc_hd__o211a_1 _20976_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_13823_),
    .C1(_14251_),
    .X(_04552_));
 sky130_fd_sc_hd__a211o_1 _20977_ (.A1(_04540_),
    .A2(\alu_shr[8] ),
    .B1(_04551_),
    .C1(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__a221o_1 _20978_ (.A1(\alu_shl[8] ),
    .A2(_04545_),
    .B1(_14797_),
    .B2(_04550_),
    .C1(_04553_),
    .X(_02142_));
 sky130_vsdinv _20979_ (.A(_14794_),
    .Y(_04554_));
 sky130_fd_sc_hd__o211a_1 _20980_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_13822_),
    .C1(_14249_),
    .X(_04555_));
 sky130_fd_sc_hd__a221o_1 _20981_ (.A1(_04554_),
    .A2(_04539_),
    .B1(_04540_),
    .B2(\alu_shr[9] ),
    .C1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__a221o_1 _20982_ (.A1(\alu_shl[9] ),
    .A2(_04545_),
    .B1(_14796_),
    .B2(_04550_),
    .C1(_04556_),
    .X(_02143_));
 sky130_fd_sc_hd__buf_4 _20983_ (.A(_04529_),
    .X(_04557_));
 sky130_fd_sc_hd__buf_4 _20984_ (.A(_04530_),
    .X(_04558_));
 sky130_fd_sc_hd__a211oi_4 _20985_ (.A1(net339),
    .A2(_14247_),
    .B1(_04557_),
    .C1(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__clkbuf_2 _20986_ (.A(_04499_),
    .X(_04560_));
 sky130_fd_sc_hd__o2bb2ai_1 _20987_ (.A1_N(_04560_),
    .A2_N(_04547_),
    .B1(_13821_),
    .B2(_14247_),
    .Y(_04561_));
 sky130_fd_sc_hd__o2bb2ai_1 _20988_ (.A1_N(\alu_shr[10] ),
    .A2_N(_04525_),
    .B1(_04559_),
    .B2(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__a221o_1 _20989_ (.A1(\alu_shl[10] ),
    .A2(_04545_),
    .B1(_14793_),
    .B2(_04550_),
    .C1(_04562_),
    .X(_02144_));
 sky130_fd_sc_hd__a211oi_4 _20990_ (.A1(_13820_),
    .A2(_14246_),
    .B1(_04557_),
    .C1(_04558_),
    .Y(_04563_));
 sky130_fd_sc_hd__o2bb2ai_1 _20991_ (.A1_N(_04560_),
    .A2_N(_04547_),
    .B1(_13820_),
    .B2(_14246_),
    .Y(_04564_));
 sky130_fd_sc_hd__o2bb2ai_1 _20992_ (.A1_N(\alu_shr[11] ),
    .A2_N(_04525_),
    .B1(_04563_),
    .B2(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__a221o_1 _20993_ (.A1(\alu_shl[11] ),
    .A2(_04545_),
    .B1(_14798_),
    .B2(_04550_),
    .C1(_04565_),
    .X(_02145_));
 sky130_fd_sc_hd__o211ai_4 _20994_ (.A1(_13007_),
    .A2(_13050_),
    .B1(_13819_),
    .C1(_14245_),
    .Y(_04566_));
 sky130_fd_sc_hd__nor3b_4 _20995_ (.A(_14808_),
    .B(_14809_),
    .C_N(_04517_),
    .Y(_04567_));
 sky130_fd_sc_hd__a221oi_2 _20996_ (.A1(\alu_shl[12] ),
    .A2(_04515_),
    .B1(_04516_),
    .B2(\alu_shr[12] ),
    .C1(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__o211ai_4 _20997_ (.A1(_14808_),
    .A2(_04501_),
    .B1(_04566_),
    .C1(_04568_),
    .Y(_02146_));
 sky130_fd_sc_hd__nor3b_2 _20998_ (.A(_14806_),
    .B(_14807_),
    .C_N(_04496_),
    .Y(_04569_));
 sky130_fd_sc_hd__a211oi_2 _20999_ (.A1(_13818_),
    .A2(_14243_),
    .B1(_13012_),
    .C1(_13053_),
    .Y(_04570_));
 sky130_fd_sc_hd__o2bb2ai_1 _21000_ (.A1_N(_04500_),
    .A2_N(_04503_),
    .B1(_13818_),
    .B2(_14243_),
    .Y(_04571_));
 sky130_fd_sc_hd__o2bb2ai_1 _21001_ (.A1_N(\alu_shr[13] ),
    .A2_N(_04516_),
    .B1(_04570_),
    .B2(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__a211o_1 _21002_ (.A1(\alu_shl[13] ),
    .A2(_04520_),
    .B1(_04569_),
    .C1(_04572_),
    .X(_02147_));
 sky130_fd_sc_hd__a211oi_4 _21003_ (.A1(_13816_),
    .A2(_14242_),
    .B1(_04557_),
    .C1(_04558_),
    .Y(_04573_));
 sky130_fd_sc_hd__o2bb2ai_1 _21004_ (.A1_N(_04560_),
    .A2_N(_04547_),
    .B1(_13816_),
    .B2(_14242_),
    .Y(_04574_));
 sky130_fd_sc_hd__o2bb2ai_1 _21005_ (.A1_N(\alu_shr[14] ),
    .A2_N(_04525_),
    .B1(_04573_),
    .B2(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__a221o_1 _21006_ (.A1(\alu_shl[14] ),
    .A2(_04545_),
    .B1(_14802_),
    .B2(_04550_),
    .C1(_04575_),
    .X(_02148_));
 sky130_fd_sc_hd__clkbuf_2 _21007_ (.A(_04514_),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_2 _21008_ (.A(_04506_),
    .X(_04577_));
 sky130_fd_sc_hd__a211oi_4 _21009_ (.A1(_13815_),
    .A2(_14241_),
    .B1(_04557_),
    .C1(_04558_),
    .Y(_04578_));
 sky130_fd_sc_hd__o2bb2ai_1 _21010_ (.A1_N(_04560_),
    .A2_N(_04547_),
    .B1(_13815_),
    .B2(_14241_),
    .Y(_04579_));
 sky130_fd_sc_hd__o2bb2ai_2 _21011_ (.A1_N(\alu_shr[15] ),
    .A2_N(_04577_),
    .B1(_04578_),
    .B2(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__a221o_1 _21012_ (.A1(\alu_shl[15] ),
    .A2(_04576_),
    .B1(_14805_),
    .B2(_04550_),
    .C1(_04580_),
    .X(_02149_));
 sky130_fd_sc_hd__clkbuf_2 _21013_ (.A(_04517_),
    .X(_04581_));
 sky130_fd_sc_hd__a211oi_2 _21014_ (.A1(_13814_),
    .A2(_14240_),
    .B1(_04557_),
    .C1(_04558_),
    .Y(_04582_));
 sky130_fd_sc_hd__o2bb2ai_1 _21015_ (.A1_N(_04560_),
    .A2_N(_04547_),
    .B1(_13814_),
    .B2(_14240_),
    .Y(_04583_));
 sky130_fd_sc_hd__o2bb2ai_1 _21016_ (.A1_N(\alu_shr[16] ),
    .A2_N(_04577_),
    .B1(_04582_),
    .B2(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__a221o_1 _21017_ (.A1(\alu_shl[16] ),
    .A2(_04576_),
    .B1(_14757_),
    .B2(_04581_),
    .C1(_04584_),
    .X(_02150_));
 sky130_fd_sc_hd__a211oi_2 _21018_ (.A1(_13813_),
    .A2(_14238_),
    .B1(_04557_),
    .C1(_04558_),
    .Y(_04585_));
 sky130_fd_sc_hd__clkbuf_2 _21019_ (.A(_04502_),
    .X(_04586_));
 sky130_fd_sc_hd__o2bb2ai_1 _21020_ (.A1_N(_04560_),
    .A2_N(_04586_),
    .B1(_13813_),
    .B2(_14238_),
    .Y(_04587_));
 sky130_fd_sc_hd__o2bb2ai_1 _21021_ (.A1_N(\alu_shr[17] ),
    .A2_N(_04577_),
    .B1(_04585_),
    .B2(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__a221o_1 _21022_ (.A1(\alu_shl[17] ),
    .A2(_04576_),
    .B1(_14756_),
    .B2(_04581_),
    .C1(_04588_),
    .X(_02151_));
 sky130_fd_sc_hd__nor2_1 _21023_ (.A(_14752_),
    .B(_14750_),
    .Y(_04589_));
 sky130_fd_sc_hd__o211a_1 _21024_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_13812_),
    .C1(_14236_),
    .X(_04590_));
 sky130_fd_sc_hd__a221o_1 _21025_ (.A1(_14753_),
    .A2(_04539_),
    .B1(_04540_),
    .B2(\alu_shr[18] ),
    .C1(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__a221o_1 _21026_ (.A1(\alu_shl[18] ),
    .A2(_04576_),
    .B1(_04589_),
    .B2(_04581_),
    .C1(_04591_),
    .X(_02152_));
 sky130_fd_sc_hd__nor2_1 _21027_ (.A(_14766_),
    .B(_14767_),
    .Y(_04592_));
 sky130_fd_sc_hd__buf_4 _21028_ (.A(_04529_),
    .X(_04593_));
 sky130_fd_sc_hd__buf_4 _21029_ (.A(_04530_),
    .X(_04594_));
 sky130_fd_sc_hd__a211oi_4 _21030_ (.A1(_13811_),
    .A2(_14234_),
    .B1(_04593_),
    .C1(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__clkbuf_2 _21031_ (.A(_04499_),
    .X(_04596_));
 sky130_fd_sc_hd__o2bb2ai_1 _21032_ (.A1_N(_04596_),
    .A2_N(_04586_),
    .B1(_13811_),
    .B2(_14234_),
    .Y(_04597_));
 sky130_fd_sc_hd__o2bb2ai_1 _21033_ (.A1_N(\alu_shr[19] ),
    .A2_N(_04577_),
    .B1(_04595_),
    .B2(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__a221o_1 _21034_ (.A1(\alu_shl[19] ),
    .A2(_04576_),
    .B1(_04592_),
    .B2(_04581_),
    .C1(_04598_),
    .X(_02153_));
 sky130_vsdinv _21035_ (.A(_14760_),
    .Y(_04599_));
 sky130_fd_sc_hd__o211a_1 _21036_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_13809_),
    .C1(_14233_),
    .X(_04600_));
 sky130_fd_sc_hd__a221o_1 _21037_ (.A1(_04599_),
    .A2(_04539_),
    .B1(_04540_),
    .B2(\alu_shr[20] ),
    .C1(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__a221o_1 _21038_ (.A1(\alu_shl[20] ),
    .A2(_04576_),
    .B1(_14762_),
    .B2(_04581_),
    .C1(_04601_),
    .X(_02154_));
 sky130_fd_sc_hd__clkbuf_2 _21039_ (.A(_04514_),
    .X(_04602_));
 sky130_fd_sc_hd__a211oi_4 _21040_ (.A1(_13808_),
    .A2(_14232_),
    .B1(_04593_),
    .C1(_04594_),
    .Y(_04603_));
 sky130_fd_sc_hd__o2bb2ai_1 _21041_ (.A1_N(_04596_),
    .A2_N(_04586_),
    .B1(_13808_),
    .B2(_14232_),
    .Y(_04604_));
 sky130_fd_sc_hd__o2bb2ai_1 _21042_ (.A1_N(\alu_shr[21] ),
    .A2_N(_04577_),
    .B1(_04603_),
    .B2(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__a221o_1 _21043_ (.A1(\alu_shl[21] ),
    .A2(_04602_),
    .B1(_14765_),
    .B2(_04581_),
    .C1(_04605_),
    .X(_02155_));
 sky130_fd_sc_hd__buf_2 _21044_ (.A(_04517_),
    .X(_04606_));
 sky130_fd_sc_hd__o22a_1 _21045_ (.A1(_04529_),
    .A2(_04530_),
    .B1(_13807_),
    .B2(_14231_),
    .X(_04607_));
 sky130_fd_sc_hd__o211a_1 _21046_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_13807_),
    .C1(_14231_),
    .X(_04608_));
 sky130_fd_sc_hd__a211o_1 _21047_ (.A1(_04540_),
    .A2(\alu_shr[22] ),
    .B1(_04607_),
    .C1(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__a221o_1 _21048_ (.A1(\alu_shl[22] ),
    .A2(_04602_),
    .B1(_14758_),
    .B2(_04606_),
    .C1(_04609_),
    .X(_02156_));
 sky130_fd_sc_hd__nor2_2 _21049_ (.A(_14768_),
    .B(_14769_),
    .Y(_04610_));
 sky130_fd_sc_hd__a211oi_2 _21050_ (.A1(_13806_),
    .A2(_14230_),
    .B1(_04593_),
    .C1(_04594_),
    .Y(_04611_));
 sky130_fd_sc_hd__o2bb2ai_1 _21051_ (.A1_N(_04596_),
    .A2_N(_04586_),
    .B1(_13806_),
    .B2(_14230_),
    .Y(_04612_));
 sky130_fd_sc_hd__o2bb2ai_1 _21052_ (.A1_N(\alu_shr[23] ),
    .A2_N(_04577_),
    .B1(_04611_),
    .B2(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__a221o_1 _21053_ (.A1(\alu_shl[23] ),
    .A2(_04602_),
    .B1(_04610_),
    .B2(_04606_),
    .C1(_04613_),
    .X(_02157_));
 sky130_fd_sc_hd__o211ai_2 _21054_ (.A1(_13007_),
    .A2(_13050_),
    .B1(_13805_),
    .C1(_14229_),
    .Y(_04614_));
 sky130_fd_sc_hd__nor3b_4 _21055_ (.A(_14727_),
    .B(_14728_),
    .C_N(_04517_),
    .Y(_04615_));
 sky130_fd_sc_hd__a221oi_2 _21056_ (.A1(\alu_shl[24] ),
    .A2(_04515_),
    .B1(_04516_),
    .B2(\alu_shr[24] ),
    .C1(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__o211ai_2 _21057_ (.A1(_14727_),
    .A2(_04501_),
    .B1(_04614_),
    .C1(_04616_),
    .Y(_02158_));
 sky130_fd_sc_hd__a211oi_4 _21058_ (.A1(_13804_),
    .A2(_14226_),
    .B1(_04593_),
    .C1(_04594_),
    .Y(_04617_));
 sky130_fd_sc_hd__o2bb2ai_1 _21059_ (.A1_N(_04596_),
    .A2_N(_04586_),
    .B1(_13804_),
    .B2(_14226_),
    .Y(_04618_));
 sky130_fd_sc_hd__o2bb2ai_1 _21060_ (.A1_N(\alu_shr[25] ),
    .A2_N(_04507_),
    .B1(_04617_),
    .B2(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__a221o_1 _21061_ (.A1(\alu_shl[25] ),
    .A2(_04602_),
    .B1(_14731_),
    .B2(_04606_),
    .C1(_04619_),
    .X(_02159_));
 sky130_fd_sc_hd__a211oi_2 _21062_ (.A1(_13801_),
    .A2(_14224_),
    .B1(_04593_),
    .C1(_04594_),
    .Y(_04620_));
 sky130_fd_sc_hd__o2bb2ai_1 _21063_ (.A1_N(_04596_),
    .A2_N(_04586_),
    .B1(_13801_),
    .B2(_14224_),
    .Y(_04621_));
 sky130_fd_sc_hd__o2bb2ai_1 _21064_ (.A1_N(\alu_shr[26] ),
    .A2_N(_04507_),
    .B1(_04620_),
    .B2(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__a221o_1 _21065_ (.A1(\alu_shl[26] ),
    .A2(_04602_),
    .B1(_14734_),
    .B2(_04606_),
    .C1(_04622_),
    .X(_02160_));
 sky130_vsdinv _21066_ (.A(_14735_),
    .Y(_04623_));
 sky130_fd_sc_hd__o211a_1 _21067_ (.A1(instr_and),
    .A2(instr_andi),
    .B1(_13800_),
    .C1(_14222_),
    .X(_04624_));
 sky130_fd_sc_hd__a221o_1 _21068_ (.A1(_04623_),
    .A2(_04539_),
    .B1(_04506_),
    .B2(\alu_shr[27] ),
    .C1(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__a221o_1 _21069_ (.A1(\alu_shl[27] ),
    .A2(_04602_),
    .B1(_14737_),
    .B2(_04606_),
    .C1(_04625_),
    .X(_02161_));
 sky130_fd_sc_hd__nor2_1 _21070_ (.A(_14741_),
    .B(_14742_),
    .Y(_04626_));
 sky130_fd_sc_hd__a211oi_4 _21071_ (.A1(_13799_),
    .A2(_14220_),
    .B1(_04593_),
    .C1(_04594_),
    .Y(_04627_));
 sky130_fd_sc_hd__o2bb2ai_1 _21072_ (.A1_N(_04596_),
    .A2_N(_04502_),
    .B1(_13799_),
    .B2(_14220_),
    .Y(_04628_));
 sky130_fd_sc_hd__o2bb2ai_1 _21073_ (.A1_N(\alu_shr[28] ),
    .A2_N(_04507_),
    .B1(_04627_),
    .B2(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__a221o_1 _21074_ (.A1(\alu_shl[28] ),
    .A2(_04515_),
    .B1(_04626_),
    .B2(_04606_),
    .C1(_04629_),
    .X(_02162_));
 sky130_fd_sc_hd__nor2_1 _21075_ (.A(_14739_),
    .B(_14740_),
    .Y(_04630_));
 sky130_fd_sc_hd__a211oi_2 _21076_ (.A1(_13798_),
    .A2(_14218_),
    .B1(_04529_),
    .C1(_04530_),
    .Y(_04631_));
 sky130_fd_sc_hd__o2bb2ai_1 _21077_ (.A1_N(_04499_),
    .A2_N(_04502_),
    .B1(_13798_),
    .B2(_14218_),
    .Y(_04632_));
 sky130_fd_sc_hd__o2bb2ai_1 _21078_ (.A1_N(\alu_shr[29] ),
    .A2_N(_04507_),
    .B1(_04631_),
    .B2(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__a221o_1 _21079_ (.A1(\alu_shl[29] ),
    .A2(_04515_),
    .B1(_04630_),
    .B2(_04496_),
    .C1(_04633_),
    .X(_02163_));
 sky130_fd_sc_hd__o211ai_1 _21080_ (.A1(_13007_),
    .A2(_13050_),
    .B1(_13797_),
    .C1(_14217_),
    .Y(_04634_));
 sky130_fd_sc_hd__nor3b_4 _21081_ (.A(_14743_),
    .B(_14744_),
    .C_N(_04495_),
    .Y(_04635_));
 sky130_fd_sc_hd__a221oi_2 _21082_ (.A1(\alu_shl[30] ),
    .A2(_04514_),
    .B1(_04516_),
    .B2(\alu_shr[30] ),
    .C1(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__o211ai_1 _21083_ (.A1(_14743_),
    .A2(_04501_),
    .B1(_04634_),
    .C1(_04636_),
    .Y(_02164_));
 sky130_fd_sc_hd__xor2_4 _21084_ (.A(net330),
    .B(_12808_),
    .X(_04637_));
 sky130_fd_sc_hd__nor2_1 _21085_ (.A(_14746_),
    .B(_04502_),
    .Y(_04638_));
 sky130_fd_sc_hd__a221o_1 _21086_ (.A1(_14745_),
    .A2(_04539_),
    .B1(_04506_),
    .B2(\alu_shr[31] ),
    .C1(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__a221o_1 _21087_ (.A1(\alu_shl[31] ),
    .A2(_04515_),
    .B1(_04637_),
    .B2(_04496_),
    .C1(_04639_),
    .X(_02165_));
 sky130_fd_sc_hd__and4_1 _21088_ (.A(_12665_),
    .B(_12636_),
    .C(_14715_),
    .D(_12631_),
    .X(_02166_));
 sky130_fd_sc_hd__buf_4 _21089_ (.A(_15157_),
    .X(_04640_));
 sky130_fd_sc_hd__a211o_4 _21090_ (.A1(_15156_),
    .A2(_04640_),
    .B1(_00304_),
    .C1(_01683_),
    .X(net233));
 sky130_fd_sc_hd__a211o_4 _21091_ (.A1(_15156_),
    .A2(_04640_),
    .B1(_01683_),
    .C1(_15160_),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 _21092_ (.A(\mem_wordsize[1] ),
    .X(_04641_));
 sky130_fd_sc_hd__buf_2 _21093_ (.A(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__a22o_1 _21094_ (.A1(_13823_),
    .A2(_04640_),
    .B1(_13840_),
    .B2(_04642_),
    .X(_02167_));
 sky130_fd_sc_hd__a22o_1 _21095_ (.A1(_13822_),
    .A2(_04640_),
    .B1(_13838_),
    .B2(_04642_),
    .X(_02168_));
 sky130_fd_sc_hd__a22o_1 _21096_ (.A1(_13821_),
    .A2(_04640_),
    .B1(_13836_),
    .B2(_04642_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _21097_ (.A1(_13820_),
    .A2(_04640_),
    .B1(_14645_),
    .B2(_04642_),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_1 _21098_ (.A1(_13819_),
    .A2(_15175_),
    .B1(_13832_),
    .B2(_04641_),
    .X(_02171_));
 sky130_fd_sc_hd__a22o_1 _21099_ (.A1(_13818_),
    .A2(_15175_),
    .B1(_13830_),
    .B2(_04641_),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_1 _21100_ (.A1(_13816_),
    .A2(_15175_),
    .B1(_13828_),
    .B2(_04641_),
    .X(_02173_));
 sky130_fd_sc_hd__a22o_1 _21101_ (.A1(_13815_),
    .A2(_15175_),
    .B1(_13826_),
    .B2(_04641_),
    .X(_02174_));
 sky130_fd_sc_hd__buf_2 _21102_ (.A(_04641_),
    .X(_04643_));
 sky130_fd_sc_hd__o21a_1 _21103_ (.A1(_04098_),
    .A2(_04643_),
    .B1(_13840_),
    .X(_02175_));
 sky130_fd_sc_hd__o21a_1 _21104_ (.A1(_04098_),
    .A2(_04643_),
    .B1(_13838_),
    .X(_02176_));
 sky130_fd_sc_hd__buf_2 _21105_ (.A(_15157_),
    .X(_04644_));
 sky130_fd_sc_hd__o21a_1 _21106_ (.A1(_04644_),
    .A2(_04643_),
    .B1(_14646_),
    .X(_02177_));
 sky130_fd_sc_hd__o21a_1 _21107_ (.A1(_04644_),
    .A2(_04643_),
    .B1(_14644_),
    .X(_02178_));
 sky130_fd_sc_hd__o21a_1 _21108_ (.A1(_04644_),
    .A2(_04643_),
    .B1(_14643_),
    .X(_02179_));
 sky130_fd_sc_hd__o21a_1 _21109_ (.A1(_04644_),
    .A2(_04643_),
    .B1(_13830_),
    .X(_02180_));
 sky130_fd_sc_hd__o21a_1 _21110_ (.A1(_04644_),
    .A2(_04642_),
    .B1(_13828_),
    .X(_02181_));
 sky130_fd_sc_hd__o21a_1 _21111_ (.A1(_04644_),
    .A2(_04642_),
    .B1(_13826_),
    .X(_02182_));
 sky130_fd_sc_hd__nand2_8 _21112_ (.A(_14837_),
    .B(_12858_),
    .Y(_02183_));
 sky130_fd_sc_hd__or2_1 _21113_ (.A(\irq_pending[3] ),
    .B(net26),
    .X(_02214_));
 sky130_fd_sc_hd__o21a_1 _21114_ (.A1(\irq_pending[3] ),
    .A2(net26),
    .B1(\irq_mask[3] ),
    .X(_02215_));
 sky130_vsdinv _21115_ (.A(_01700_),
    .Y(_02217_));
 sky130_fd_sc_hd__or2_1 _21116_ (.A(\irq_pending[4] ),
    .B(net27),
    .X(_02218_));
 sky130_fd_sc_hd__o21a_1 _21117_ (.A1(\irq_pending[4] ),
    .A2(net27),
    .B1(\irq_mask[4] ),
    .X(_02219_));
 sky130_fd_sc_hd__or2_1 _21118_ (.A(\irq_pending[5] ),
    .B(net28),
    .X(_02221_));
 sky130_fd_sc_hd__o21a_1 _21119_ (.A1(\irq_pending[5] ),
    .A2(net28),
    .B1(\irq_mask[5] ),
    .X(_02222_));
 sky130_fd_sc_hd__or2_1 _21120_ (.A(\irq_pending[6] ),
    .B(net29),
    .X(_02224_));
 sky130_fd_sc_hd__o21a_1 _21121_ (.A1(\irq_pending[6] ),
    .A2(net29),
    .B1(\irq_mask[6] ),
    .X(_02225_));
 sky130_fd_sc_hd__or2_1 _21122_ (.A(\irq_pending[7] ),
    .B(net501),
    .X(_02227_));
 sky130_fd_sc_hd__o21a_1 _21123_ (.A1(\irq_pending[7] ),
    .A2(net501),
    .B1(\irq_mask[7] ),
    .X(_02228_));
 sky130_fd_sc_hd__or2_1 _21124_ (.A(\irq_pending[8] ),
    .B(net31),
    .X(_02230_));
 sky130_fd_sc_hd__o21a_1 _21125_ (.A1(\irq_pending[8] ),
    .A2(net31),
    .B1(\irq_mask[8] ),
    .X(_02231_));
 sky130_fd_sc_hd__or2_1 _21126_ (.A(\irq_pending[9] ),
    .B(net32),
    .X(_02233_));
 sky130_fd_sc_hd__o21a_1 _21127_ (.A1(\irq_pending[9] ),
    .A2(net32),
    .B1(\irq_mask[9] ),
    .X(_02234_));
 sky130_fd_sc_hd__or2_1 _21128_ (.A(\irq_pending[10] ),
    .B(net504),
    .X(_02236_));
 sky130_fd_sc_hd__o21a_1 _21129_ (.A1(\irq_pending[10] ),
    .A2(net504),
    .B1(\irq_mask[10] ),
    .X(_02237_));
 sky130_fd_sc_hd__or2_1 _21130_ (.A(\irq_pending[11] ),
    .B(net3),
    .X(_02239_));
 sky130_fd_sc_hd__o21a_1 _21131_ (.A1(\irq_pending[11] ),
    .A2(net3),
    .B1(\irq_mask[11] ),
    .X(_02240_));
 sky130_fd_sc_hd__or2_1 _21132_ (.A(\irq_pending[12] ),
    .B(net4),
    .X(_02242_));
 sky130_fd_sc_hd__o21a_1 _21133_ (.A1(\irq_pending[12] ),
    .A2(net4),
    .B1(\irq_mask[12] ),
    .X(_02243_));
 sky130_fd_sc_hd__or2_1 _21134_ (.A(\irq_pending[13] ),
    .B(net5),
    .X(_02245_));
 sky130_fd_sc_hd__o21a_1 _21135_ (.A1(\irq_pending[13] ),
    .A2(net5),
    .B1(\irq_mask[13] ),
    .X(_02246_));
 sky130_fd_sc_hd__or2_1 _21136_ (.A(\irq_pending[14] ),
    .B(net6),
    .X(_02248_));
 sky130_fd_sc_hd__o21a_1 _21137_ (.A1(\irq_pending[14] ),
    .A2(net6),
    .B1(\irq_mask[14] ),
    .X(_02249_));
 sky130_fd_sc_hd__or2_1 _21138_ (.A(\irq_pending[15] ),
    .B(net496),
    .X(_02251_));
 sky130_fd_sc_hd__o21a_1 _21139_ (.A1(\irq_pending[15] ),
    .A2(net496),
    .B1(\irq_mask[15] ),
    .X(_02252_));
 sky130_fd_sc_hd__or2_1 _21140_ (.A(\irq_pending[16] ),
    .B(net8),
    .X(_02254_));
 sky130_fd_sc_hd__o21a_1 _21141_ (.A1(\irq_pending[16] ),
    .A2(net8),
    .B1(\irq_mask[16] ),
    .X(_02255_));
 sky130_fd_sc_hd__or2_1 _21142_ (.A(\irq_pending[17] ),
    .B(net9),
    .X(_02257_));
 sky130_fd_sc_hd__o21a_1 _21143_ (.A1(\irq_pending[17] ),
    .A2(net9),
    .B1(\irq_mask[17] ),
    .X(_02258_));
 sky130_fd_sc_hd__or2_1 _21144_ (.A(\irq_pending[18] ),
    .B(net10),
    .X(_02260_));
 sky130_fd_sc_hd__o21a_1 _21145_ (.A1(\irq_pending[18] ),
    .A2(net10),
    .B1(\irq_mask[18] ),
    .X(_02261_));
 sky130_fd_sc_hd__or2_1 _21146_ (.A(\irq_pending[19] ),
    .B(net11),
    .X(_02263_));
 sky130_fd_sc_hd__o21a_1 _21147_ (.A1(\irq_pending[19] ),
    .A2(net11),
    .B1(\irq_mask[19] ),
    .X(_02264_));
 sky130_fd_sc_hd__or2_1 _21148_ (.A(\irq_pending[20] ),
    .B(net505),
    .X(_02266_));
 sky130_fd_sc_hd__o21a_1 _21149_ (.A1(\irq_pending[20] ),
    .A2(net505),
    .B1(\irq_mask[20] ),
    .X(_02267_));
 sky130_fd_sc_hd__or2_1 _21150_ (.A(\irq_pending[21] ),
    .B(net14),
    .X(_02269_));
 sky130_fd_sc_hd__o21a_1 _21151_ (.A1(\irq_pending[21] ),
    .A2(net14),
    .B1(\irq_mask[21] ),
    .X(_02270_));
 sky130_fd_sc_hd__or2_1 _21152_ (.A(\irq_pending[22] ),
    .B(net15),
    .X(_02272_));
 sky130_fd_sc_hd__o21a_1 _21153_ (.A1(\irq_pending[22] ),
    .A2(net15),
    .B1(\irq_mask[22] ),
    .X(_02273_));
 sky130_fd_sc_hd__or2_1 _21154_ (.A(\irq_pending[23] ),
    .B(net16),
    .X(_02275_));
 sky130_fd_sc_hd__o21a_1 _21155_ (.A1(\irq_pending[23] ),
    .A2(net16),
    .B1(\irq_mask[23] ),
    .X(_02276_));
 sky130_fd_sc_hd__or2_1 _21156_ (.A(\irq_pending[24] ),
    .B(net17),
    .X(_02278_));
 sky130_fd_sc_hd__o21a_1 _21157_ (.A1(\irq_pending[24] ),
    .A2(net17),
    .B1(\irq_mask[24] ),
    .X(_02279_));
 sky130_fd_sc_hd__or2_1 _21158_ (.A(\irq_pending[25] ),
    .B(net18),
    .X(_02281_));
 sky130_fd_sc_hd__o21a_1 _21159_ (.A1(\irq_pending[25] ),
    .A2(net18),
    .B1(\irq_mask[25] ),
    .X(_02282_));
 sky130_fd_sc_hd__or2_1 _21160_ (.A(\irq_pending[26] ),
    .B(net19),
    .X(_02284_));
 sky130_fd_sc_hd__o21a_1 _21161_ (.A1(\irq_pending[26] ),
    .A2(net19),
    .B1(\irq_mask[26] ),
    .X(_02285_));
 sky130_fd_sc_hd__or2_1 _21162_ (.A(\irq_pending[27] ),
    .B(net503),
    .X(_02287_));
 sky130_fd_sc_hd__o21a_1 _21163_ (.A1(\irq_pending[27] ),
    .A2(net503),
    .B1(\irq_mask[27] ),
    .X(_02288_));
 sky130_fd_sc_hd__or2_1 _21164_ (.A(\irq_pending[28] ),
    .B(net502),
    .X(_02290_));
 sky130_fd_sc_hd__o21a_1 _21165_ (.A1(\irq_pending[28] ),
    .A2(net502),
    .B1(\irq_mask[28] ),
    .X(_02291_));
 sky130_fd_sc_hd__or2_1 _21166_ (.A(\irq_pending[29] ),
    .B(net22),
    .X(_02293_));
 sky130_fd_sc_hd__o21a_1 _21167_ (.A1(\irq_pending[29] ),
    .A2(net22),
    .B1(\irq_mask[29] ),
    .X(_02294_));
 sky130_fd_sc_hd__or2_1 _21168_ (.A(\irq_pending[30] ),
    .B(net24),
    .X(_02296_));
 sky130_fd_sc_hd__o21a_1 _21169_ (.A1(\irq_pending[30] ),
    .A2(net24),
    .B1(\irq_mask[30] ),
    .X(_02297_));
 sky130_fd_sc_hd__or2_1 _21170_ (.A(\irq_pending[31] ),
    .B(net25),
    .X(_02299_));
 sky130_fd_sc_hd__o21a_1 _21171_ (.A1(\irq_pending[31] ),
    .A2(net25),
    .B1(\irq_mask[31] ),
    .X(_02300_));
 sky130_fd_sc_hd__nor3_1 _21172_ (.A(_14843_),
    .B(_14838_),
    .C(_14841_),
    .Y(_04645_));
 sky130_fd_sc_hd__and3b_1 _21173_ (.A_N(_14842_),
    .B(_14857_),
    .C(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__nor3b_2 _21174_ (.A(\timer[1] ),
    .B(_14844_),
    .C_N(\timer[0] ),
    .Y(_04647_));
 sky130_fd_sc_hd__and4b_1 _21175_ (.A_N(\timer[6] ),
    .B(_14846_),
    .C(_14847_),
    .D(_14850_),
    .X(_04648_));
 sky130_fd_sc_hd__and4_1 _21176_ (.A(_04647_),
    .B(_14852_),
    .C(_04648_),
    .D(_14855_),
    .X(_04649_));
 sky130_fd_sc_hd__a21o_1 _21177_ (.A1(_04646_),
    .A2(_04649_),
    .B1(\irq_pending[0] ),
    .X(_02302_));
 sky130_fd_sc_hd__or2_1 _21178_ (.A(_02303_),
    .B(net1),
    .X(_02304_));
 sky130_fd_sc_hd__o21a_1 _21179_ (.A1(_02303_),
    .A2(net1),
    .B1(\irq_mask[0] ),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_1 _21180_ (.A(\irq_pending[2] ),
    .B(net23),
    .Y(_02307_));
 sky130_fd_sc_hd__o21ai_1 _21181_ (.A1(\irq_pending[2] ),
    .A2(net23),
    .B1(_13537_),
    .Y(_02308_));
 sky130_fd_sc_hd__nor2b_1 _21182_ (.A(_02310_),
    .B_N(_12650_),
    .Y(_02311_));
 sky130_fd_sc_hd__o22ai_1 _21183_ (.A1(_14651_),
    .A2(_13537_),
    .B1(_02310_),
    .B2(_13322_),
    .Y(_02312_));
 sky130_fd_sc_hd__o21bai_1 _21184_ (.A1(_14651_),
    .A2(_13537_),
    .B1_N(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__o21bai_1 _21185_ (.A1(_14651_),
    .A2(_13537_),
    .B1_N(_02316_),
    .Y(_02317_));
 sky130_vsdinv _21186_ (.A(_12808_),
    .Y(_04650_));
 sky130_fd_sc_hd__inv_2 _21187_ (.A(_13797_),
    .Y(_02405_));
 sky130_fd_sc_hd__and2b_1 _21188_ (.A_N(_14219_),
    .B(net358),
    .X(_04651_));
 sky130_fd_sc_hd__and2b_1 _21189_ (.A_N(_14223_),
    .B(net356),
    .X(_04652_));
 sky130_fd_sc_hd__and2b_1 _21190_ (.A_N(_14228_),
    .B(net354),
    .X(_04653_));
 sky130_fd_sc_hd__o21ai_1 _21191_ (.A1(_14729_),
    .A2(_14730_),
    .B1(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__or2b_1 _21192_ (.A(_14225_),
    .B_N(net355),
    .X(_04655_));
 sky130_fd_sc_hd__a21oi_1 _21193_ (.A1(_04654_),
    .A2(_04655_),
    .B1(_14734_),
    .Y(_04656_));
 sky130_fd_sc_hd__o21bai_1 _21194_ (.A1(_04652_),
    .A2(_04656_),
    .B1_N(_14737_),
    .Y(_04657_));
 sky130_fd_sc_hd__or2b_1 _21195_ (.A(_14222_),
    .B_N(_13800_),
    .X(_04658_));
 sky130_fd_sc_hd__a21oi_1 _21196_ (.A1(_04657_),
    .A2(_04658_),
    .B1(_04626_),
    .Y(_04659_));
 sky130_fd_sc_hd__o21bai_1 _21197_ (.A1(_04651_),
    .A2(_04659_),
    .B1_N(_04630_),
    .Y(_04660_));
 sky130_fd_sc_hd__nand2_1 _21198_ (.A(_15000_),
    .B(net359),
    .Y(_04661_));
 sky130_fd_sc_hd__a21bo_1 _21199_ (.A1(_04660_),
    .A2(_04661_),
    .B1_N(_14747_),
    .X(_04662_));
 sky130_fd_sc_hd__o31a_1 _21200_ (.A1(_02405_),
    .A2(net329),
    .A3(_04637_),
    .B1(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__and2b_1 _21201_ (.A_N(_14233_),
    .B(_13809_),
    .X(_04664_));
 sky130_fd_sc_hd__and2b_1 _21202_ (.A_N(_14236_),
    .B(_13812_),
    .X(_04665_));
 sky130_fd_sc_hd__and2b_1 _21203_ (.A_N(_14239_),
    .B(net345),
    .X(_04666_));
 sky130_fd_sc_hd__o21ai_1 _21204_ (.A1(_14754_),
    .A2(_14755_),
    .B1(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__or2b_1 _21205_ (.A(_14238_),
    .B_N(net346),
    .X(_04668_));
 sky130_fd_sc_hd__a21oi_1 _21206_ (.A1(_04667_),
    .A2(_04668_),
    .B1(_04589_),
    .Y(_04669_));
 sky130_fd_sc_hd__o21bai_1 _21207_ (.A1(_04665_),
    .A2(_04669_),
    .B1_N(_04592_),
    .Y(_04670_));
 sky130_fd_sc_hd__or2b_1 _21208_ (.A(_14234_),
    .B_N(_13811_),
    .X(_04671_));
 sky130_fd_sc_hd__a21oi_1 _21209_ (.A1(_04670_),
    .A2(_04671_),
    .B1(_14762_),
    .Y(_04672_));
 sky130_fd_sc_hd__o21bai_1 _21210_ (.A1(_04664_),
    .A2(_04672_),
    .B1_N(_14765_),
    .Y(_04673_));
 sky130_fd_sc_hd__or2b_1 _21211_ (.A(_14232_),
    .B_N(net351),
    .X(_04674_));
 sky130_fd_sc_hd__a21o_1 _21212_ (.A1(_04673_),
    .A2(_04674_),
    .B1(_14758_),
    .X(_04675_));
 sky130_fd_sc_hd__or2b_1 _21213_ (.A(_14231_),
    .B_N(_13807_),
    .X(_04676_));
 sky130_fd_sc_hd__a21oi_2 _21214_ (.A1(_04675_),
    .A2(_04676_),
    .B1(_04610_),
    .Y(_04677_));
 sky130_fd_sc_hd__and2b_1 _21215_ (.A_N(_14230_),
    .B(_13806_),
    .X(_04678_));
 sky130_fd_sc_hd__and2b_1 _21216_ (.A_N(_14241_),
    .B(net344),
    .X(_04679_));
 sky130_fd_sc_hd__inv_2 _21217_ (.A(net342),
    .Y(_02354_));
 sky130_fd_sc_hd__inv_2 _21218_ (.A(_13819_),
    .Y(_02351_));
 sky130_fd_sc_hd__o21bai_1 _21219_ (.A1(_14806_),
    .A2(_14807_),
    .B1_N(_14245_),
    .Y(_04680_));
 sky130_fd_sc_hd__o22ai_1 _21220_ (.A1(_02354_),
    .A2(_14243_),
    .B1(_02351_),
    .B2(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__o21ai_1 _21221_ (.A1(_14800_),
    .A2(_14801_),
    .B1(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__or2b_1 _21222_ (.A(_14242_),
    .B_N(net343),
    .X(_04683_));
 sky130_fd_sc_hd__a21oi_1 _21223_ (.A1(_04682_),
    .A2(_04683_),
    .B1(_14805_),
    .Y(_04684_));
 sky130_fd_sc_hd__and2b_1 _21224_ (.A_N(_14250_),
    .B(net368),
    .X(_04685_));
 sky130_fd_sc_hd__o21ai_1 _21225_ (.A1(_14794_),
    .A2(_14795_),
    .B1(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__or2b_1 _21226_ (.A(_14249_),
    .B_N(net369),
    .X(_04687_));
 sky130_fd_sc_hd__a21o_1 _21227_ (.A1(_04686_),
    .A2(_04687_),
    .B1(_14793_),
    .X(_04688_));
 sky130_fd_sc_hd__or2b_1 _21228_ (.A(_14247_),
    .B_N(net339),
    .X(_04689_));
 sky130_fd_sc_hd__a21oi_1 _21229_ (.A1(_04688_),
    .A2(_04689_),
    .B1(_14798_),
    .Y(_04690_));
 sky130_fd_sc_hd__and2b_1 _21230_ (.A_N(_14246_),
    .B(net340),
    .X(_04691_));
 sky130_fd_sc_hd__and2b_1 _21231_ (.A_N(_14256_),
    .B(_13827_),
    .X(_04692_));
 sky130_fd_sc_hd__and2b_1 _21232_ (.A_N(_14258_),
    .B(_13831_),
    .X(_04693_));
 sky130_fd_sc_hd__and2b_1 _21233_ (.A_N(_14260_),
    .B(_13833_),
    .X(_04694_));
 sky130_fd_sc_hd__o21a_1 _21234_ (.A1(_02318_),
    .A2(_00048_),
    .B1(net317),
    .X(_04695_));
 sky130_fd_sc_hd__or2b_1 _21235_ (.A(_14261_),
    .B_N(_13835_),
    .X(_04696_));
 sky130_fd_sc_hd__o31ai_1 _21236_ (.A1(_00049_),
    .A2(_14787_),
    .A3(_04695_),
    .B1(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__o21a_1 _21237_ (.A1(_14779_),
    .A2(_14780_),
    .B1(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__o21ba_1 _21238_ (.A1(_04694_),
    .A2(_04698_),
    .B1_N(_14791_),
    .X(_04699_));
 sky130_fd_sc_hd__o21bai_1 _21239_ (.A1(_04693_),
    .A2(_04699_),
    .B1_N(_04534_),
    .Y(_04700_));
 sky130_fd_sc_hd__or2b_1 _21240_ (.A(_14257_),
    .B_N(_13829_),
    .X(_04701_));
 sky130_fd_sc_hd__a21oi_1 _21241_ (.A1(_04700_),
    .A2(_04701_),
    .B1(_14790_),
    .Y(_04702_));
 sky130_fd_sc_hd__o21bai_1 _21242_ (.A1(_04692_),
    .A2(_04702_),
    .B1_N(_14786_),
    .Y(_04703_));
 sky130_fd_sc_hd__or2b_1 _21243_ (.A(_14253_),
    .B_N(_13825_),
    .X(_04704_));
 sky130_fd_sc_hd__a21oi_1 _21244_ (.A1(_04703_),
    .A2(_04704_),
    .B1(_14799_),
    .Y(_04705_));
 sky130_fd_sc_hd__o31a_1 _21245_ (.A1(_04690_),
    .A2(_04691_),
    .A3(_04705_),
    .B1(_14811_),
    .X(_04706_));
 sky130_fd_sc_hd__o311a_1 _21246_ (.A1(_04679_),
    .A2(_04684_),
    .A3(_04706_),
    .B1(_14759_),
    .C1(_14771_),
    .X(_04707_));
 sky130_fd_sc_hd__o31ai_4 _21247_ (.A1(_04677_),
    .A2(_04678_),
    .A3(_04707_),
    .B1(_14749_),
    .Y(_04708_));
 sky130_fd_sc_hd__o211a_1 _21248_ (.A1(_12797_),
    .A2(_04650_),
    .B1(_04663_),
    .C1(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__nor2_1 _21249_ (.A(_00000_),
    .B(_04709_),
    .Y(_00002_));
 sky130_vsdinv _21250_ (.A(_00000_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand3b_1 _21251_ (.A_N(_04637_),
    .B(_04708_),
    .C(_04663_),
    .Y(_04711_));
 sky130_fd_sc_hd__o211a_1 _21252_ (.A1(_12797_),
    .A2(_04650_),
    .B1(_04710_),
    .C1(_04711_),
    .X(_00001_));
 sky130_fd_sc_hd__buf_2 _21253_ (.A(\pcpi_mul.rs2[0] ),
    .X(_04712_));
 sky130_fd_sc_hd__buf_2 _21254_ (.A(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__buf_6 _21255_ (.A(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__buf_6 _21256_ (.A(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__buf_4 _21257_ (.A(\pcpi_mul.rs1[0] ),
    .X(_04716_));
 sky130_fd_sc_hd__buf_4 _21258_ (.A(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__buf_4 _21259_ (.A(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__buf_6 _21260_ (.A(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__clkbuf_4 _21261_ (.A(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__buf_2 _21262_ (.A(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__and2_1 _21263_ (.A(_04715_),
    .B(_04721_),
    .X(_02623_));
 sky130_fd_sc_hd__xnor2_1 _21264_ (.A(_13837_),
    .B(_13839_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _21265_ (.A(_15170_),
    .B(net200),
    .Y(_04722_));
 sky130_fd_sc_hd__xor2_2 _21266_ (.A(net317),
    .B(_02320_),
    .X(_04723_));
 sky130_fd_sc_hd__xor2_1 _21267_ (.A(_04722_),
    .B(_04723_),
    .X(_02602_));
 sky130_fd_sc_hd__nor2_4 _21268_ (.A(net491),
    .B(net200),
    .Y(_04724_));
 sky130_fd_sc_hd__xor2_1 _21269_ (.A(_13836_),
    .B(_04724_),
    .X(_02322_));
 sky130_fd_sc_hd__xor2_1 _21270_ (.A(_14262_),
    .B(_02323_),
    .X(_04725_));
 sky130_fd_sc_hd__and2_1 _21271_ (.A(net317),
    .B(_02320_),
    .X(_04726_));
 sky130_fd_sc_hd__a21o_1 _21272_ (.A1(_04723_),
    .A2(_04722_),
    .B1(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__xor2_1 _21273_ (.A(_04725_),
    .B(_04727_),
    .X(_02613_));
 sky130_fd_sc_hd__nor3_4 _21274_ (.A(_13835_),
    .B(_13837_),
    .C(_13839_),
    .Y(_04728_));
 sky130_fd_sc_hd__xor2_1 _21275_ (.A(_13834_),
    .B(_04728_),
    .X(_02325_));
 sky130_fd_sc_hd__nor2_1 _21276_ (.A(net331),
    .B(_02326_),
    .Y(_04729_));
 sky130_fd_sc_hd__and2_1 _21277_ (.A(net331),
    .B(_02326_),
    .X(_04730_));
 sky130_fd_sc_hd__nor2_1 _21278_ (.A(_04729_),
    .B(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__or2_1 _21279_ (.A(net328),
    .B(_02323_),
    .X(_04732_));
 sky130_fd_sc_hd__and2_1 _21280_ (.A(_14261_),
    .B(_02323_),
    .X(_04733_));
 sky130_fd_sc_hd__a21o_1 _21281_ (.A1(_04727_),
    .A2(_04732_),
    .B1(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__xor2_1 _21282_ (.A(_04731_),
    .B(_04734_),
    .X(_02616_));
 sky130_fd_sc_hd__nand3_4 _21283_ (.A(_04724_),
    .B(_14648_),
    .C(_14649_),
    .Y(_04735_));
 sky130_fd_sc_hd__xor2_1 _21284_ (.A(_02327_),
    .B(_04735_),
    .X(_02328_));
 sky130_fd_sc_hd__xor2_1 _21285_ (.A(_14259_),
    .B(_02329_),
    .X(_04736_));
 sky130_vsdinv _21286_ (.A(_04729_),
    .Y(_04737_));
 sky130_fd_sc_hd__a21o_1 _21287_ (.A1(_04734_),
    .A2(_04737_),
    .B1(_04730_),
    .X(_04738_));
 sky130_fd_sc_hd__xor2_1 _21288_ (.A(_04736_),
    .B(_04738_),
    .X(_02617_));
 sky130_fd_sc_hd__inv_2 _21289_ (.A(_13830_),
    .Y(_02330_));
 sky130_fd_sc_hd__nand3_4 _21290_ (.A(_04728_),
    .B(_14647_),
    .C(_14648_),
    .Y(_04739_));
 sky130_fd_sc_hd__xor2_1 _21291_ (.A(_02330_),
    .B(_04739_),
    .X(_02331_));
 sky130_fd_sc_hd__nor2_1 _21292_ (.A(net333),
    .B(_02332_),
    .Y(_04740_));
 sky130_fd_sc_hd__and2_1 _21293_ (.A(net333),
    .B(_02332_),
    .X(_04741_));
 sky130_fd_sc_hd__nor2_1 _21294_ (.A(_04740_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__or2_1 _21295_ (.A(net332),
    .B(_02329_),
    .X(_04743_));
 sky130_fd_sc_hd__and2_1 _21296_ (.A(_14258_),
    .B(_02329_),
    .X(_04744_));
 sky130_fd_sc_hd__a21o_1 _21297_ (.A1(_04738_),
    .A2(_04743_),
    .B1(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__xor2_1 _21298_ (.A(_04742_),
    .B(_04745_),
    .X(_02618_));
 sky130_fd_sc_hd__inv_2 _21299_ (.A(net228),
    .Y(_02333_));
 sky130_fd_sc_hd__nor3_4 _21300_ (.A(net227),
    .B(net226),
    .C(_04735_),
    .Y(_04746_));
 sky130_fd_sc_hd__xor2_1 _21301_ (.A(_13828_),
    .B(_04746_),
    .X(_02334_));
 sky130_fd_sc_hd__xor2_2 _21302_ (.A(net334),
    .B(_02335_),
    .X(_04747_));
 sky130_vsdinv _21303_ (.A(_04740_),
    .Y(_04748_));
 sky130_fd_sc_hd__a21o_1 _21304_ (.A1(_04745_),
    .A2(_04748_),
    .B1(_04741_),
    .X(_04749_));
 sky130_fd_sc_hd__xor2_1 _21305_ (.A(_04747_),
    .B(_04749_),
    .X(_02619_));
 sky130_fd_sc_hd__inv_2 _21306_ (.A(net229),
    .Y(_02336_));
 sky130_fd_sc_hd__nor3_4 _21307_ (.A(_13827_),
    .B(_13829_),
    .C(_04739_),
    .Y(_04750_));
 sky130_fd_sc_hd__xor2_1 _21308_ (.A(_13826_),
    .B(_04750_),
    .X(_02337_));
 sky130_fd_sc_hd__xnor2_1 _21309_ (.A(net335),
    .B(_02338_),
    .Y(_04751_));
 sky130_fd_sc_hd__and2_1 _21310_ (.A(_14256_),
    .B(_02335_),
    .X(_04752_));
 sky130_fd_sc_hd__a21oi_1 _21311_ (.A1(_04749_),
    .A2(_04747_),
    .B1(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__xor2_1 _21312_ (.A(_04751_),
    .B(_04753_),
    .X(_02620_));
 sky130_fd_sc_hd__inv_2 _21313_ (.A(_13823_),
    .Y(_02339_));
 sky130_fd_sc_hd__nand3_4 _21314_ (.A(_04746_),
    .B(_02336_),
    .C(_02333_),
    .Y(_04754_));
 sky130_fd_sc_hd__xor2_1 _21315_ (.A(_02339_),
    .B(_04754_),
    .X(_02340_));
 sky130_fd_sc_hd__xor2_2 _21316_ (.A(net336),
    .B(_02341_),
    .X(_04755_));
 sky130_fd_sc_hd__and2b_1 _21317_ (.A_N(_04751_),
    .B(_04747_),
    .X(_04756_));
 sky130_fd_sc_hd__o211a_1 _21318_ (.A1(_14252_),
    .A2(_02338_),
    .B1(_14255_),
    .C1(_02335_),
    .X(_04757_));
 sky130_fd_sc_hd__a221oi_2 _21319_ (.A1(_14252_),
    .A2(_02338_),
    .B1(_04749_),
    .B2(_04756_),
    .C1(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__xnor2_1 _21320_ (.A(_04755_),
    .B(_04758_),
    .Y(_02621_));
 sky130_fd_sc_hd__inv_2 _21321_ (.A(_13822_),
    .Y(_02342_));
 sky130_fd_sc_hd__nand3_4 _21322_ (.A(_04750_),
    .B(_02339_),
    .C(_02336_),
    .Y(_04759_));
 sky130_fd_sc_hd__xor2_1 _21323_ (.A(_02342_),
    .B(_04759_),
    .X(_02343_));
 sky130_fd_sc_hd__xnor2_2 _21324_ (.A(net337),
    .B(_02344_),
    .Y(_04760_));
 sky130_fd_sc_hd__and2b_1 _21325_ (.A_N(_04758_),
    .B(_04755_),
    .X(_04761_));
 sky130_fd_sc_hd__a21oi_1 _21326_ (.A1(_14251_),
    .A2(_02341_),
    .B1(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__xor2_1 _21327_ (.A(_04760_),
    .B(_04762_),
    .X(_02622_));
 sky130_fd_sc_hd__inv_2 _21328_ (.A(net339),
    .Y(_02345_));
 sky130_fd_sc_hd__nor3_4 _21329_ (.A(net369),
    .B(net368),
    .C(_04754_),
    .Y(_04763_));
 sky130_fd_sc_hd__xor2_1 _21330_ (.A(_13821_),
    .B(_04763_),
    .X(_02346_));
 sky130_fd_sc_hd__xor2_2 _21331_ (.A(net307),
    .B(_02347_),
    .X(_04764_));
 sky130_fd_sc_hd__o211a_1 _21332_ (.A1(_14248_),
    .A2(_02344_),
    .B1(_14250_),
    .C1(_02341_),
    .X(_04765_));
 sky130_fd_sc_hd__nor3b_2 _21333_ (.A(_04760_),
    .B(_04758_),
    .C_N(_04755_),
    .Y(_04766_));
 sky130_fd_sc_hd__a211o_1 _21334_ (.A1(_14248_),
    .A2(_02344_),
    .B1(_04765_),
    .C1(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__xor2_1 _21335_ (.A(_04764_),
    .B(_04767_),
    .X(_02592_));
 sky130_fd_sc_hd__inv_2 _21336_ (.A(net340),
    .Y(_02348_));
 sky130_fd_sc_hd__nor3_2 _21337_ (.A(_13821_),
    .B(_13822_),
    .C(_04759_),
    .Y(_04768_));
 sky130_fd_sc_hd__xor2_1 _21338_ (.A(_13820_),
    .B(_04768_),
    .X(_02349_));
 sky130_fd_sc_hd__xor2_2 _21339_ (.A(net308),
    .B(_02350_),
    .X(_04769_));
 sky130_fd_sc_hd__and2_1 _21340_ (.A(net307),
    .B(_02347_),
    .X(_04770_));
 sky130_fd_sc_hd__a21o_1 _21341_ (.A1(_04767_),
    .A2(_04764_),
    .B1(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__xor2_1 _21342_ (.A(_04769_),
    .B(_04771_),
    .X(_02593_));
 sky130_fd_sc_hd__nand3_4 _21343_ (.A(_04763_),
    .B(_02348_),
    .C(_02345_),
    .Y(_04772_));
 sky130_fd_sc_hd__xor2_1 _21344_ (.A(_02351_),
    .B(_04772_),
    .X(_02352_));
 sky130_fd_sc_hd__xor2_2 _21345_ (.A(net309),
    .B(_02353_),
    .X(_04773_));
 sky130_fd_sc_hd__and2_1 _21346_ (.A(net308),
    .B(_02350_),
    .X(_04774_));
 sky130_fd_sc_hd__a21o_1 _21347_ (.A1(_04771_),
    .A2(_04769_),
    .B1(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__xor2_1 _21348_ (.A(_04773_),
    .B(_04775_),
    .X(_02594_));
 sky130_fd_sc_hd__nor2_2 _21349_ (.A(_13819_),
    .B(_04772_),
    .Y(_04776_));
 sky130_fd_sc_hd__xor2_1 _21350_ (.A(_13818_),
    .B(_04776_),
    .X(_02355_));
 sky130_fd_sc_hd__xor2_2 _21351_ (.A(net310),
    .B(_02356_),
    .X(_04777_));
 sky130_fd_sc_hd__and2_1 _21352_ (.A(_04775_),
    .B(_04773_),
    .X(_04778_));
 sky130_fd_sc_hd__a21o_1 _21353_ (.A1(net309),
    .A2(_02353_),
    .B1(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__xor2_1 _21354_ (.A(_04777_),
    .B(_04779_),
    .X(_02595_));
 sky130_fd_sc_hd__inv_2 _21355_ (.A(net343),
    .Y(_02357_));
 sky130_fd_sc_hd__nor3_4 _21356_ (.A(net342),
    .B(net341),
    .C(_04772_),
    .Y(_04780_));
 sky130_fd_sc_hd__xor2_1 _21357_ (.A(_13816_),
    .B(_04780_),
    .X(_02358_));
 sky130_fd_sc_hd__nor2_2 _21358_ (.A(net311),
    .B(_02359_),
    .Y(_04781_));
 sky130_fd_sc_hd__and2_2 _21359_ (.A(net311),
    .B(_02359_),
    .X(_04782_));
 sky130_fd_sc_hd__nor2_4 _21360_ (.A(_04781_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__and2_1 _21361_ (.A(net310),
    .B(_02356_),
    .X(_04784_));
 sky130_fd_sc_hd__a21o_1 _21362_ (.A1(_04779_),
    .A2(_04777_),
    .B1(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__xor2_1 _21363_ (.A(_04783_),
    .B(_04785_),
    .X(_02596_));
 sky130_fd_sc_hd__inv_2 _21364_ (.A(net344),
    .Y(_02360_));
 sky130_fd_sc_hd__and3_1 _21365_ (.A(_04776_),
    .B(_02357_),
    .C(_02354_),
    .X(_04786_));
 sky130_fd_sc_hd__xor2_1 _21366_ (.A(_13815_),
    .B(_04786_),
    .X(_02361_));
 sky130_fd_sc_hd__xnor2_2 _21367_ (.A(net312),
    .B(_02362_),
    .Y(_04787_));
 sky130_fd_sc_hd__a21oi_4 _21368_ (.A1(_04785_),
    .A2(_04783_),
    .B1(_04782_),
    .Y(_04788_));
 sky130_fd_sc_hd__xor2_1 _21369_ (.A(_04787_),
    .B(_04788_),
    .X(_02597_));
 sky130_fd_sc_hd__inv_2 _21370_ (.A(_13814_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand3_4 _21371_ (.A(_04780_),
    .B(_02360_),
    .C(_02357_),
    .Y(_04789_));
 sky130_fd_sc_hd__xor2_1 _21372_ (.A(_02363_),
    .B(_04789_),
    .X(_02364_));
 sky130_fd_sc_hd__xor2_2 _21373_ (.A(_14239_),
    .B(_02365_),
    .X(_04790_));
 sky130_fd_sc_hd__and2_1 _21374_ (.A(net312),
    .B(_02362_),
    .X(_04791_));
 sky130_fd_sc_hd__o21bai_4 _21375_ (.A1(_04787_),
    .A2(_04788_),
    .B1_N(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__xor2_1 _21376_ (.A(_04790_),
    .B(_04792_),
    .X(_02598_));
 sky130_vsdinv _21377_ (.A(_13813_),
    .Y(_02366_));
 sky130_fd_sc_hd__nor2_1 _21378_ (.A(_13814_),
    .B(_04789_),
    .Y(_04793_));
 sky130_fd_sc_hd__xor2_1 _21379_ (.A(_13813_),
    .B(_04793_),
    .X(_02367_));
 sky130_fd_sc_hd__xnor2_1 _21380_ (.A(net314),
    .B(_02368_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand2_1 _21381_ (.A(_04792_),
    .B(_04790_),
    .Y(_04795_));
 sky130_fd_sc_hd__a21boi_1 _21382_ (.A1(_14240_),
    .A2(_02365_),
    .B1_N(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__xor2_1 _21383_ (.A(_04794_),
    .B(_04796_),
    .X(_02599_));
 sky130_fd_sc_hd__inv_2 _21384_ (.A(net347),
    .Y(_02369_));
 sky130_fd_sc_hd__nor3_4 _21385_ (.A(net346),
    .B(net345),
    .C(_04789_),
    .Y(_04797_));
 sky130_fd_sc_hd__xor2_1 _21386_ (.A(_13812_),
    .B(_04797_),
    .X(_02370_));
 sky130_fd_sc_hd__xnor2_2 _21387_ (.A(net315),
    .B(_02371_),
    .Y(_04798_));
 sky130_fd_sc_hd__and2b_1 _21388_ (.A_N(_04794_),
    .B(_04790_),
    .X(_04799_));
 sky130_fd_sc_hd__and2_1 _21389_ (.A(_14237_),
    .B(_02368_),
    .X(_04800_));
 sky130_fd_sc_hd__o211a_1 _21390_ (.A1(_14237_),
    .A2(_02368_),
    .B1(_14239_),
    .C1(_02365_),
    .X(_04801_));
 sky130_fd_sc_hd__a211oi_4 _21391_ (.A1(_04792_),
    .A2(_04799_),
    .B1(_04800_),
    .C1(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__xor2_1 _21392_ (.A(_04798_),
    .B(_04802_),
    .X(_02600_));
 sky130_fd_sc_hd__inv_2 _21393_ (.A(net348),
    .Y(_02372_));
 sky130_fd_sc_hd__and4_1 _21394_ (.A(_04776_),
    .B(_02360_),
    .C(_02357_),
    .D(_02354_),
    .X(_04803_));
 sky130_fd_sc_hd__and4_1 _21395_ (.A(_04803_),
    .B(_02369_),
    .C(_02366_),
    .D(_02363_),
    .X(_04804_));
 sky130_fd_sc_hd__xor2_1 _21396_ (.A(_13811_),
    .B(_04804_),
    .X(_02373_));
 sky130_fd_sc_hd__nor2_1 _21397_ (.A(net316),
    .B(_02374_),
    .Y(_04805_));
 sky130_fd_sc_hd__and2_1 _21398_ (.A(net316),
    .B(_02374_),
    .X(_04806_));
 sky130_fd_sc_hd__nor2_2 _21399_ (.A(_04805_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__and2_1 _21400_ (.A(net315),
    .B(_02371_),
    .X(_04808_));
 sky130_fd_sc_hd__o21bai_2 _21401_ (.A1(_04798_),
    .A2(_04802_),
    .B1_N(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__xor2_1 _21402_ (.A(_04807_),
    .B(_04809_),
    .X(_02601_));
 sky130_fd_sc_hd__inv_2 _21403_ (.A(_13809_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand3_4 _21404_ (.A(_04797_),
    .B(_02372_),
    .C(_02369_),
    .Y(_04810_));
 sky130_fd_sc_hd__xor2_1 _21405_ (.A(_02375_),
    .B(_04810_),
    .X(_02376_));
 sky130_fd_sc_hd__xnor2_2 _21406_ (.A(net318),
    .B(_02377_),
    .Y(_04811_));
 sky130_fd_sc_hd__a21oi_2 _21407_ (.A1(_04809_),
    .A2(_04807_),
    .B1(_04806_),
    .Y(_04812_));
 sky130_fd_sc_hd__xor2_1 _21408_ (.A(_04811_),
    .B(_04812_),
    .X(_02603_));
 sky130_vsdinv _21409_ (.A(_13808_),
    .Y(_02378_));
 sky130_fd_sc_hd__nor2_1 _21410_ (.A(_13809_),
    .B(_04810_),
    .Y(_04813_));
 sky130_fd_sc_hd__xor2_1 _21411_ (.A(_13808_),
    .B(_04813_),
    .X(_02379_));
 sky130_fd_sc_hd__nor2_1 _21412_ (.A(net319),
    .B(_02380_),
    .Y(_04814_));
 sky130_fd_sc_hd__and2_1 _21413_ (.A(net319),
    .B(_02380_),
    .X(_04815_));
 sky130_fd_sc_hd__nor2_2 _21414_ (.A(_04814_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__and2_1 _21415_ (.A(net318),
    .B(_02377_),
    .X(_04817_));
 sky130_fd_sc_hd__o21bai_2 _21416_ (.A1(_04811_),
    .A2(_04812_),
    .B1_N(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__xor2_1 _21417_ (.A(_04816_),
    .B(_04818_),
    .X(_02604_));
 sky130_fd_sc_hd__inv_2 _21418_ (.A(net352),
    .Y(_02381_));
 sky130_fd_sc_hd__nor3_4 _21419_ (.A(net351),
    .B(net350),
    .C(_04810_),
    .Y(_04819_));
 sky130_fd_sc_hd__xor2_1 _21420_ (.A(_13807_),
    .B(_04819_),
    .X(_02382_));
 sky130_fd_sc_hd__xnor2_1 _21421_ (.A(net320),
    .B(_02383_),
    .Y(_04820_));
 sky130_fd_sc_hd__a21oi_2 _21422_ (.A1(_04818_),
    .A2(_04816_),
    .B1(_04815_),
    .Y(_04821_));
 sky130_fd_sc_hd__xor2_1 _21423_ (.A(_04820_),
    .B(_04821_),
    .X(_02605_));
 sky130_fd_sc_hd__inv_2 _21424_ (.A(net353),
    .Y(_02384_));
 sky130_fd_sc_hd__and4_1 _21425_ (.A(_04793_),
    .B(_02372_),
    .C(_02369_),
    .D(_02366_),
    .X(_04822_));
 sky130_fd_sc_hd__and4_1 _21426_ (.A(_04822_),
    .B(_02381_),
    .C(_02378_),
    .D(_02375_),
    .X(_04823_));
 sky130_fd_sc_hd__xor2_1 _21427_ (.A(_13806_),
    .B(_04823_),
    .X(_02385_));
 sky130_fd_sc_hd__nor2_2 _21428_ (.A(net321),
    .B(_02386_),
    .Y(_04824_));
 sky130_fd_sc_hd__and2_2 _21429_ (.A(net321),
    .B(_02386_),
    .X(_04825_));
 sky130_fd_sc_hd__nor2_4 _21430_ (.A(_04824_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__and2_1 _21431_ (.A(net320),
    .B(_02383_),
    .X(_04827_));
 sky130_fd_sc_hd__o21bai_2 _21432_ (.A1(_04820_),
    .A2(_04821_),
    .B1_N(_04827_),
    .Y(_04828_));
 sky130_fd_sc_hd__xor2_1 _21433_ (.A(_04826_),
    .B(_04828_),
    .X(_02606_));
 sky130_fd_sc_hd__inv_2 _21434_ (.A(_13805_),
    .Y(_02387_));
 sky130_fd_sc_hd__nand3_4 _21435_ (.A(_04819_),
    .B(_02384_),
    .C(_02381_),
    .Y(_04829_));
 sky130_fd_sc_hd__xor2_1 _21436_ (.A(_02387_),
    .B(_04829_),
    .X(_02388_));
 sky130_fd_sc_hd__xor2_2 _21437_ (.A(_14228_),
    .B(_02389_),
    .X(_04830_));
 sky130_fd_sc_hd__a21oi_4 _21438_ (.A1(_04828_),
    .A2(_04826_),
    .B1(_04825_),
    .Y(_04831_));
 sky130_fd_sc_hd__xnor2_1 _21439_ (.A(_04830_),
    .B(_04831_),
    .Y(_02607_));
 sky130_fd_sc_hd__inv_2 _21440_ (.A(_13804_),
    .Y(_02390_));
 sky130_fd_sc_hd__nor2_2 _21441_ (.A(_13805_),
    .B(_04829_),
    .Y(_04832_));
 sky130_fd_sc_hd__xor2_1 _21442_ (.A(_13804_),
    .B(_04832_),
    .X(_02391_));
 sky130_fd_sc_hd__xor2_2 _21443_ (.A(_14225_),
    .B(_02392_),
    .X(_04833_));
 sky130_fd_sc_hd__and2b_1 _21444_ (.A_N(_04831_),
    .B(_04830_),
    .X(_04834_));
 sky130_fd_sc_hd__a21oi_1 _21445_ (.A1(_14229_),
    .A2(_02389_),
    .B1(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__xnor2_1 _21446_ (.A(_04833_),
    .B(_04835_),
    .Y(_02608_));
 sky130_fd_sc_hd__inv_2 _21447_ (.A(_13801_),
    .Y(_02393_));
 sky130_fd_sc_hd__nor3_4 _21448_ (.A(net355),
    .B(_13805_),
    .C(_04829_),
    .Y(_04836_));
 sky130_fd_sc_hd__xor2_1 _21449_ (.A(_13801_),
    .B(_04836_),
    .X(_02394_));
 sky130_fd_sc_hd__xor2_4 _21450_ (.A(_14223_),
    .B(_02395_),
    .X(_04837_));
 sky130_fd_sc_hd__nand2_1 _21451_ (.A(_04830_),
    .B(_04833_),
    .Y(_04838_));
 sky130_fd_sc_hd__o211a_1 _21452_ (.A1(net323),
    .A2(_02392_),
    .B1(net322),
    .C1(_02389_),
    .X(_04839_));
 sky130_fd_sc_hd__a21o_1 _21453_ (.A1(_14226_),
    .A2(_02392_),
    .B1(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__o21bai_4 _21454_ (.A1(_04838_),
    .A2(_04831_),
    .B1_N(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__xor2_1 _21455_ (.A(_04837_),
    .B(_04841_),
    .X(_02609_));
 sky130_fd_sc_hd__inv_2 _21456_ (.A(_13800_),
    .Y(_02396_));
 sky130_fd_sc_hd__nand3_1 _21457_ (.A(_04832_),
    .B(_02393_),
    .C(_02390_),
    .Y(_04842_));
 sky130_fd_sc_hd__xor2_1 _21458_ (.A(_02396_),
    .B(_04842_),
    .X(_02397_));
 sky130_fd_sc_hd__xnor2_1 _21459_ (.A(_14221_),
    .B(_02398_),
    .Y(_04843_));
 sky130_fd_sc_hd__and2_1 _21460_ (.A(_14224_),
    .B(_02395_),
    .X(_04844_));
 sky130_fd_sc_hd__a21oi_1 _21461_ (.A1(_04841_),
    .A2(_04837_),
    .B1(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__xor2_1 _21462_ (.A(_04843_),
    .B(_04845_),
    .X(_02610_));
 sky130_fd_sc_hd__inv_2 _21463_ (.A(_13799_),
    .Y(_02399_));
 sky130_fd_sc_hd__nand3_4 _21464_ (.A(_04836_),
    .B(_02396_),
    .C(_02393_),
    .Y(_04846_));
 sky130_fd_sc_hd__xor2_1 _21465_ (.A(_02399_),
    .B(_04846_),
    .X(_02400_));
 sky130_fd_sc_hd__xnor2_1 _21466_ (.A(_14220_),
    .B(_02401_),
    .Y(_04847_));
 sky130_fd_sc_hd__and2b_1 _21467_ (.A_N(_04843_),
    .B(_04837_),
    .X(_04848_));
 sky130_fd_sc_hd__o211a_1 _21468_ (.A1(_14221_),
    .A2(_02398_),
    .B1(_14223_),
    .C1(_02395_),
    .X(_04849_));
 sky130_fd_sc_hd__a21oi_1 _21469_ (.A1(_14222_),
    .A2(_02398_),
    .B1(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__a21boi_4 _21470_ (.A1(_04841_),
    .A2(_04848_),
    .B1_N(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__xor2_1 _21471_ (.A(_04847_),
    .B(_04851_),
    .X(_02611_));
 sky130_fd_sc_hd__inv_2 _21472_ (.A(net359),
    .Y(_02402_));
 sky130_fd_sc_hd__nor2_1 _21473_ (.A(net358),
    .B(_04846_),
    .Y(_04852_));
 sky130_fd_sc_hd__xor2_1 _21474_ (.A(_13798_),
    .B(_04852_),
    .X(_02403_));
 sky130_fd_sc_hd__nor2_1 _21475_ (.A(net327),
    .B(_02404_),
    .Y(_04853_));
 sky130_fd_sc_hd__and2_1 _21476_ (.A(net327),
    .B(_02404_),
    .X(_04854_));
 sky130_fd_sc_hd__nor2_1 _21477_ (.A(_04853_),
    .B(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__nor2_2 _21478_ (.A(_14219_),
    .B(_02401_),
    .Y(_04856_));
 sky130_fd_sc_hd__and2_1 _21479_ (.A(_14219_),
    .B(_02401_),
    .X(_04857_));
 sky130_fd_sc_hd__o21bai_4 _21480_ (.A1(_04856_),
    .A2(_04851_),
    .B1_N(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__xor2_1 _21481_ (.A(_04855_),
    .B(_04858_),
    .X(_02612_));
 sky130_fd_sc_hd__nor3_2 _21482_ (.A(_13798_),
    .B(_13799_),
    .C(_04846_),
    .Y(_04859_));
 sky130_fd_sc_hd__xor2_1 _21483_ (.A(_13797_),
    .B(_04859_),
    .X(_02406_));
 sky130_fd_sc_hd__xnor2_1 _21484_ (.A(_14217_),
    .B(_02407_),
    .Y(_04860_));
 sky130_vsdinv _21485_ (.A(_04853_),
    .Y(_04861_));
 sky130_fd_sc_hd__a21oi_4 _21486_ (.A1(_04858_),
    .A2(_04861_),
    .B1(_04854_),
    .Y(_04862_));
 sky130_fd_sc_hd__xor2_1 _21487_ (.A(_04860_),
    .B(_04862_),
    .X(_02614_));
 sky130_fd_sc_hd__nand3_1 _21488_ (.A(_04852_),
    .B(_02405_),
    .C(_02402_),
    .Y(_04863_));
 sky130_fd_sc_hd__xor2_1 _21489_ (.A(_12808_),
    .B(_04863_),
    .X(_02408_));
 sky130_fd_sc_hd__nor2_1 _21490_ (.A(_14217_),
    .B(_02407_),
    .Y(_04864_));
 sky130_fd_sc_hd__and2_1 _21491_ (.A(net329),
    .B(_02407_),
    .X(_04865_));
 sky130_fd_sc_hd__o21bai_1 _21492_ (.A1(_04864_),
    .A2(_04862_),
    .B1_N(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__xnor2_1 _21493_ (.A(_12797_),
    .B(_02409_),
    .Y(_04867_));
 sky130_vsdinv _21494_ (.A(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand2_1 _21495_ (.A(_04866_),
    .B(_04868_),
    .Y(_04869_));
 sky130_vsdinv _21496_ (.A(_04865_),
    .Y(_04870_));
 sky130_fd_sc_hd__o211ai_1 _21497_ (.A1(_04864_),
    .A2(_04862_),
    .B1(_04870_),
    .C1(_04867_),
    .Y(_04871_));
 sky130_fd_sc_hd__nand2_1 _21498_ (.A(_04869_),
    .B(_04871_),
    .Y(_02615_));
 sky130_fd_sc_hd__buf_4 _21499_ (.A(_14448_),
    .X(_04872_));
 sky130_fd_sc_hd__buf_6 _21500_ (.A(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__buf_2 _21501_ (.A(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_2 _21502_ (.A(_04715_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__clkbuf_4 _21503_ (.A(_14093_),
    .X(_04876_));
 sky130_fd_sc_hd__buf_4 _21504_ (.A(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__buf_6 _21505_ (.A(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__buf_6 _21506_ (.A(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__buf_8 _21507_ (.A(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__nand2_2 _21508_ (.A(_04880_),
    .B(_04721_),
    .Y(_04881_));
 sky130_fd_sc_hd__xor2_2 _21509_ (.A(_04875_),
    .B(_04881_),
    .X(_02624_));
 sky130_fd_sc_hd__nor2_2 _21510_ (.A(_04875_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__nand2_1 _21511_ (.A(_04878_),
    .B(_04874_),
    .Y(_04883_));
 sky130_fd_sc_hd__clkbuf_4 _21512_ (.A(\pcpi_mul.rs2[2] ),
    .X(_04884_));
 sky130_fd_sc_hd__buf_4 _21513_ (.A(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__buf_6 _21514_ (.A(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__nand2_1 _21515_ (.A(_04886_),
    .B(_04719_),
    .Y(_04887_));
 sky130_fd_sc_hd__xnor2_1 _21516_ (.A(_04883_),
    .B(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__clkbuf_4 _21517_ (.A(_14441_),
    .X(_04889_));
 sky130_fd_sc_hd__clkbuf_4 _21518_ (.A(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__buf_4 _21519_ (.A(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__nand3b_4 _21520_ (.A_N(_04888_),
    .B(_04715_),
    .C(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__o21ai_1 _21521_ (.A1(_14098_),
    .A2(_14445_),
    .B1(_04888_),
    .Y(_04893_));
 sky130_fd_sc_hd__and2_1 _21522_ (.A(_04892_),
    .B(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__xor2_1 _21523_ (.A(_04882_),
    .B(_04894_),
    .X(_02625_));
 sky130_fd_sc_hd__nand3_2 _21524_ (.A(_04892_),
    .B(_04882_),
    .C(_04893_),
    .Y(_04895_));
 sky130_fd_sc_hd__nor2_2 _21525_ (.A(_04883_),
    .B(_04887_),
    .Y(_04896_));
 sky130_fd_sc_hd__clkbuf_4 _21526_ (.A(\pcpi_mul.rs1[3] ),
    .X(_04897_));
 sky130_fd_sc_hd__buf_2 _21527_ (.A(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__buf_2 _21528_ (.A(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__buf_4 _21529_ (.A(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__and2_2 _21530_ (.A(_04715_),
    .B(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__nand2_4 _21531_ (.A(_14084_),
    .B(_04718_),
    .Y(_04902_));
 sky130_fd_sc_hd__nand3_4 _21532_ (.A(_04885_),
    .B(_04877_),
    .C(_04873_),
    .Y(_04903_));
 sky130_fd_sc_hd__buf_4 _21533_ (.A(\pcpi_mul.rs2[2] ),
    .X(_04904_));
 sky130_fd_sc_hd__buf_4 _21534_ (.A(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__clkbuf_4 _21535_ (.A(\pcpi_mul.rs1[1] ),
    .X(_04906_));
 sky130_fd_sc_hd__buf_4 _21536_ (.A(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__buf_6 _21537_ (.A(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__buf_4 _21538_ (.A(\pcpi_mul.rs2[1] ),
    .X(_04909_));
 sky130_fd_sc_hd__buf_4 _21539_ (.A(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__a22o_1 _21540_ (.A1(_04905_),
    .A2(_04908_),
    .B1(_04910_),
    .B2(_04891_),
    .X(_04911_));
 sky130_fd_sc_hd__o21ai_4 _21541_ (.A1(_14444_),
    .A2(_04903_),
    .B1(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__xnor2_4 _21542_ (.A(_04902_),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__xor2_4 _21543_ (.A(_04901_),
    .B(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__xor2_1 _21544_ (.A(_04892_),
    .B(_04914_),
    .X(_04915_));
 sky130_vsdinv _21545_ (.A(_04896_),
    .Y(_04916_));
 sky130_fd_sc_hd__nor2_1 _21546_ (.A(_04916_),
    .B(_04914_),
    .Y(_04917_));
 sky130_fd_sc_hd__o21bai_2 _21547_ (.A1(_04896_),
    .A2(_04915_),
    .B1_N(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__xor2_1 _21548_ (.A(_04895_),
    .B(_04918_),
    .X(_02626_));
 sky130_fd_sc_hd__nor2_2 _21549_ (.A(_04895_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__a21o_2 _21550_ (.A1(_04916_),
    .A2(_04892_),
    .B1(_04914_),
    .X(_04920_));
 sky130_fd_sc_hd__o22ai_4 _21551_ (.A1(_14445_),
    .A2(_04903_),
    .B1(_04902_),
    .B2(_04912_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand3b_4 _21552_ (.A_N(_04913_),
    .B(_04715_),
    .C(_04900_),
    .Y(_04922_));
 sky130_fd_sc_hd__buf_4 _21553_ (.A(\pcpi_mul.rs2[4] ),
    .X(_04923_));
 sky130_fd_sc_hd__buf_4 _21554_ (.A(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__nand2_4 _21555_ (.A(_04924_),
    .B(_04716_),
    .Y(_04925_));
 sky130_fd_sc_hd__buf_2 _21556_ (.A(\pcpi_mul.rs1[4] ),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_4 _21557_ (.A(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__buf_6 _21558_ (.A(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__buf_4 _21559_ (.A(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__nand2_2 _21560_ (.A(_04714_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__xnor2_4 _21561_ (.A(_04925_),
    .B(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__buf_2 _21562_ (.A(\pcpi_mul.rs2[3] ),
    .X(_04932_));
 sky130_fd_sc_hd__clkbuf_2 _21563_ (.A(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__nand2_2 _21564_ (.A(_04933_),
    .B(_04873_),
    .Y(_04934_));
 sky130_fd_sc_hd__or4_4 _21565_ (.A(_14091_),
    .B(_14094_),
    .C(_14438_),
    .D(_14443_),
    .X(_04935_));
 sky130_fd_sc_hd__buf_4 _21566_ (.A(_14090_),
    .X(_04936_));
 sky130_fd_sc_hd__buf_4 _21567_ (.A(_04890_),
    .X(_04937_));
 sky130_fd_sc_hd__buf_4 _21568_ (.A(_14093_),
    .X(_04938_));
 sky130_fd_sc_hd__a22o_1 _21569_ (.A1(_04936_),
    .A2(_04937_),
    .B1(_04938_),
    .B2(_04899_),
    .X(_04939_));
 sky130_fd_sc_hd__nand2_2 _21570_ (.A(_04935_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__xnor2_4 _21571_ (.A(_04934_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__xnor2_4 _21572_ (.A(_04931_),
    .B(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__xor2_4 _21573_ (.A(_04922_),
    .B(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__xnor2_4 _21574_ (.A(_04921_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__xor2_4 _21575_ (.A(_04920_),
    .B(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__xor2_1 _21576_ (.A(_04919_),
    .B(_04945_),
    .X(_02627_));
 sky130_fd_sc_hd__buf_6 _21577_ (.A(_04886_),
    .X(_04946_));
 sky130_fd_sc_hd__buf_6 _21578_ (.A(_04878_),
    .X(_04947_));
 sky130_fd_sc_hd__clkbuf_4 _21579_ (.A(\pcpi_mul.rs1[3] ),
    .X(_04948_));
 sky130_fd_sc_hd__buf_4 _21580_ (.A(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__nand2_2 _21581_ (.A(\pcpi_mul.rs2[2] ),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__nand2_2 _21582_ (.A(\pcpi_mul.rs2[1] ),
    .B(_04927_),
    .Y(_04951_));
 sky130_fd_sc_hd__xnor2_4 _21583_ (.A(_04950_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__nor3_4 _21584_ (.A(_14085_),
    .B(_14445_),
    .C(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__a41oi_4 _21585_ (.A1(_04946_),
    .A2(_04947_),
    .A3(_04929_),
    .A4(_04900_),
    .B1(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__buf_4 _21586_ (.A(_04712_),
    .X(_04955_));
 sky130_fd_sc_hd__buf_4 _21587_ (.A(_04926_),
    .X(_04956_));
 sky130_fd_sc_hd__buf_4 _21588_ (.A(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__nand3b_4 _21589_ (.A_N(_04925_),
    .B(_04955_),
    .C(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__clkbuf_2 _21590_ (.A(\pcpi_mul.rs1[5] ),
    .X(_04959_));
 sky130_fd_sc_hd__buf_4 _21591_ (.A(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__nand2_2 _21592_ (.A(_04712_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__buf_2 _21593_ (.A(\pcpi_mul.rs2[5] ),
    .X(_04962_));
 sky130_fd_sc_hd__nand3_4 _21594_ (.A(_04962_),
    .B(_04923_),
    .C(_14447_),
    .Y(_04963_));
 sky130_fd_sc_hd__a22o_1 _21595_ (.A1(\pcpi_mul.rs2[5] ),
    .A2(\pcpi_mul.rs1[0] ),
    .B1(\pcpi_mul.rs2[4] ),
    .B2(_14447_),
    .X(_04964_));
 sky130_fd_sc_hd__o21ai_4 _21596_ (.A1(_14451_),
    .A2(_04963_),
    .B1(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__xnor2_4 _21597_ (.A(_04961_),
    .B(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__xnor2_4 _21598_ (.A(_04958_),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__clkbuf_4 _21599_ (.A(_14441_),
    .X(_04968_));
 sky130_fd_sc_hd__buf_2 _21600_ (.A(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__and2_2 _21601_ (.A(\pcpi_mul.rs2[3] ),
    .B(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__xnor2_4 _21602_ (.A(_04970_),
    .B(_04952_),
    .Y(_04971_));
 sky130_fd_sc_hd__or2b_1 _21603_ (.A(_04967_),
    .B_N(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__o21ai_2 _21604_ (.A1(_04958_),
    .A2(_04966_),
    .B1(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__buf_4 _21605_ (.A(_04949_),
    .X(_04974_));
 sky130_fd_sc_hd__and2_2 _21606_ (.A(_14082_),
    .B(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__clkbuf_4 _21607_ (.A(_04956_),
    .X(_04976_));
 sky130_fd_sc_hd__nand2_2 _21608_ (.A(_14090_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__buf_4 _21609_ (.A(_14426_),
    .X(_04978_));
 sky130_fd_sc_hd__nand2_2 _21610_ (.A(_14093_),
    .B(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__xnor2_4 _21611_ (.A(_04977_),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__xor2_4 _21612_ (.A(_04975_),
    .B(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__o22a_2 _21613_ (.A1(_14452_),
    .A2(_04963_),
    .B1(_04961_),
    .B2(_04965_),
    .X(_04982_));
 sky130_fd_sc_hd__clkbuf_4 _21614_ (.A(_14420_),
    .X(_04983_));
 sky130_fd_sc_hd__and2_2 _21615_ (.A(_04712_),
    .B(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__clkbuf_4 _21616_ (.A(\pcpi_mul.rs2[5] ),
    .X(_04985_));
 sky130_fd_sc_hd__buf_4 _21617_ (.A(\pcpi_mul.rs1[1] ),
    .X(_04986_));
 sky130_fd_sc_hd__nand2_2 _21618_ (.A(_04985_),
    .B(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__buf_2 _21619_ (.A(\pcpi_mul.rs1[2] ),
    .X(_04988_));
 sky130_fd_sc_hd__nand2_2 _21620_ (.A(_04923_),
    .B(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__xnor2_4 _21621_ (.A(_04987_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__xor2_4 _21622_ (.A(_04984_),
    .B(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__xnor2_4 _21623_ (.A(_04982_),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__xor2_2 _21624_ (.A(_04981_),
    .B(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__xnor2_1 _21625_ (.A(_04973_),
    .B(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__nor2_1 _21626_ (.A(_04954_),
    .B(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__buf_4 _21627_ (.A(\pcpi_mul.rs2[6] ),
    .X(_04996_));
 sky130_fd_sc_hd__buf_4 _21628_ (.A(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__buf_6 _21629_ (.A(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__buf_6 _21630_ (.A(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__and2_1 _21631_ (.A(_04999_),
    .B(_04720_),
    .X(_05000_));
 sky130_fd_sc_hd__nand2_1 _21632_ (.A(_04994_),
    .B(_04954_),
    .Y(_05001_));
 sky130_fd_sc_hd__and3b_2 _21633_ (.A_N(_04995_),
    .B(_05000_),
    .C(_05001_),
    .X(_05002_));
 sky130_vsdinv _21634_ (.A(_04995_),
    .Y(_05003_));
 sky130_fd_sc_hd__a21o_1 _21635_ (.A1(_05003_),
    .A2(_05001_),
    .B1(_05000_),
    .X(_05004_));
 sky130_fd_sc_hd__o21a_2 _21636_ (.A1(_04934_),
    .A2(_04940_),
    .B1(_04935_),
    .X(_05005_));
 sky130_fd_sc_hd__or2_4 _21637_ (.A(_04931_),
    .B(_04941_),
    .X(_05006_));
 sky130_fd_sc_hd__xnor2_4 _21638_ (.A(_04971_),
    .B(_04967_),
    .Y(_05007_));
 sky130_fd_sc_hd__xor2_4 _21639_ (.A(_05006_),
    .B(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__and2b_1 _21640_ (.A_N(_05006_),
    .B(_05007_),
    .X(_05009_));
 sky130_fd_sc_hd__o21bai_2 _21641_ (.A1(_05005_),
    .A2(_05008_),
    .B1_N(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__and3b_1 _21642_ (.A_N(_05002_),
    .B(_05004_),
    .C(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__clkbuf_2 _21643_ (.A(_05011_),
    .X(_05012_));
 sky130_vsdinv _21644_ (.A(_05002_),
    .Y(_05013_));
 sky130_fd_sc_hd__a21oi_4 _21645_ (.A1(_05013_),
    .A2(_05004_),
    .B1(_05010_),
    .Y(_05014_));
 sky130_vsdinv _21646_ (.A(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__nor2_1 _21647_ (.A(_04922_),
    .B(_04942_),
    .Y(_05016_));
 sky130_fd_sc_hd__a21o_1 _21648_ (.A1(_04943_),
    .A2(_04921_),
    .B1(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__xor2_4 _21649_ (.A(_05005_),
    .B(_05008_),
    .X(_05018_));
 sky130_fd_sc_hd__or2_1 _21650_ (.A(_05017_),
    .B(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__nor2_1 _21651_ (.A(_04920_),
    .B(_04944_),
    .Y(_05020_));
 sky130_fd_sc_hd__and2_1 _21652_ (.A(_05018_),
    .B(_05017_),
    .X(_05021_));
 sky130_fd_sc_hd__a21oi_1 _21653_ (.A1(_05019_),
    .A2(_05020_),
    .B1(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand3b_1 _21654_ (.A_N(_05012_),
    .B(_05015_),
    .C(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__o21bai_1 _21655_ (.A1(_05014_),
    .A2(_05012_),
    .B1_N(_05022_),
    .Y(_05024_));
 sky130_fd_sc_hd__xnor2_2 _21656_ (.A(_05017_),
    .B(_05018_),
    .Y(_05025_));
 sky130_fd_sc_hd__nand3b_1 _21657_ (.A_N(_05025_),
    .B(_04919_),
    .C(_04945_),
    .Y(_05026_));
 sky130_fd_sc_hd__a21oi_1 _21658_ (.A1(_05023_),
    .A2(_05024_),
    .B1(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__and3_1 _21659_ (.A(_05023_),
    .B(_05026_),
    .C(_05024_),
    .X(_05028_));
 sky130_fd_sc_hd__nor2_1 _21660_ (.A(_05027_),
    .B(_05028_),
    .Y(_02683_));
 sky130_fd_sc_hd__nor2_1 _21661_ (.A(_05014_),
    .B(_05012_),
    .Y(_05029_));
 sky130_fd_sc_hd__nor3_2 _21662_ (.A(_04944_),
    .B(_04920_),
    .C(_05025_),
    .Y(_05030_));
 sky130_fd_sc_hd__a21o_1 _21663_ (.A1(_05029_),
    .A2(_05030_),
    .B1(_05027_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_4 _21664_ (.A(_04960_),
    .X(_05032_));
 sky130_fd_sc_hd__buf_4 _21665_ (.A(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__nor3_4 _21666_ (.A(_14086_),
    .B(_14439_),
    .C(_04980_),
    .Y(_05034_));
 sky130_fd_sc_hd__a41oi_4 _21667_ (.A1(_04946_),
    .A2(_04879_),
    .A3(_05033_),
    .A4(_04929_),
    .B1(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__nor2_1 _21668_ (.A(_04982_),
    .B(_04991_),
    .Y(_05036_));
 sky130_fd_sc_hd__o21bai_4 _21669_ (.A1(_04981_),
    .A2(_04992_),
    .B1_N(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__and2_2 _21670_ (.A(_04932_),
    .B(_04928_),
    .X(_05038_));
 sky130_fd_sc_hd__buf_4 _21671_ (.A(_04978_),
    .X(_05039_));
 sky130_fd_sc_hd__nand2_2 _21672_ (.A(_04904_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__buf_4 _21673_ (.A(_04983_),
    .X(_05041_));
 sky130_fd_sc_hd__nand2_2 _21674_ (.A(_04909_),
    .B(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__xnor2_4 _21675_ (.A(_05040_),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__xor2_4 _21676_ (.A(_05038_),
    .B(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__buf_4 _21677_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05045_));
 sky130_fd_sc_hd__buf_2 _21678_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05046_));
 sky130_fd_sc_hd__buf_2 _21679_ (.A(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__buf_4 _21680_ (.A(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__and2_2 _21681_ (.A(_05045_),
    .B(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__buf_4 _21682_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05050_));
 sky130_fd_sc_hd__buf_4 _21683_ (.A(\pcpi_mul.rs1[3] ),
    .X(_05051_));
 sky130_fd_sc_hd__nand2_2 _21684_ (.A(_05050_),
    .B(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__and2_1 _21685_ (.A(_04962_),
    .B(_04988_),
    .X(_05053_));
 sky130_fd_sc_hd__xor2_4 _21686_ (.A(_05052_),
    .B(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__xor2_4 _21687_ (.A(_05049_),
    .B(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_4 _21688_ (.A(_14096_),
    .X(_05056_));
 sky130_fd_sc_hd__buf_4 _21689_ (.A(_14421_),
    .X(_05057_));
 sky130_fd_sc_hd__o32a_4 _21690_ (.A1(_05056_),
    .A2(_05057_),
    .A3(_04990_),
    .B1(_14444_),
    .B2(_04963_),
    .X(_05058_));
 sky130_fd_sc_hd__xnor2_4 _21691_ (.A(_05055_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__xor2_4 _21692_ (.A(_05044_),
    .B(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__xnor2_2 _21693_ (.A(_05037_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__nor2_4 _21694_ (.A(_05035_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__buf_4 _21695_ (.A(_14065_),
    .X(_05063_));
 sky130_fd_sc_hd__buf_6 _21696_ (.A(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__buf_6 _21697_ (.A(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__nand2_2 _21698_ (.A(_05065_),
    .B(_04718_),
    .Y(_05066_));
 sky130_fd_sc_hd__nand2_2 _21699_ (.A(_04999_),
    .B(_04874_),
    .Y(_05067_));
 sky130_fd_sc_hd__xor2_1 _21700_ (.A(_05066_),
    .B(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_1 _21701_ (.A(_05061_),
    .B(_05035_),
    .Y(_05069_));
 sky130_fd_sc_hd__and3b_2 _21702_ (.A_N(_05062_),
    .B(_05068_),
    .C(_05069_),
    .X(_05070_));
 sky130_vsdinv _21703_ (.A(_05070_),
    .Y(_05071_));
 sky130_vsdinv _21704_ (.A(_05062_),
    .Y(_05072_));
 sky130_fd_sc_hd__a21o_1 _21705_ (.A1(_05072_),
    .A2(_05069_),
    .B1(_05068_),
    .X(_05073_));
 sky130_fd_sc_hd__a21oi_1 _21706_ (.A1(_05071_),
    .A2(_05073_),
    .B1(_05002_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand3b_4 _21707_ (.A_N(_05070_),
    .B(_05073_),
    .C(_05002_),
    .Y(_05075_));
 sky130_vsdinv _21708_ (.A(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__nand2_1 _21709_ (.A(_04993_),
    .B(_04973_),
    .Y(_05077_));
 sky130_fd_sc_hd__o21a_1 _21710_ (.A1(_04954_),
    .A2(_04994_),
    .B1(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__o21a_2 _21711_ (.A1(_05074_),
    .A2(_05076_),
    .B1(_05078_),
    .X(_05079_));
 sky130_vsdinv _21712_ (.A(_05078_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand3b_4 _21713_ (.A_N(_05074_),
    .B(_05075_),
    .C(_05080_),
    .Y(_05081_));
 sky130_vsdinv _21714_ (.A(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__a21oi_1 _21715_ (.A1(_05015_),
    .A2(_05021_),
    .B1(_05012_),
    .Y(_05083_));
 sky130_fd_sc_hd__o21bai_1 _21716_ (.A1(_05079_),
    .A2(_05082_),
    .B1_N(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__nand3b_1 _21717_ (.A_N(_05079_),
    .B(_05081_),
    .C(_05083_),
    .Y(_05085_));
 sky130_fd_sc_hd__nand2_1 _21718_ (.A(_05084_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__xor2_1 _21719_ (.A(_05031_),
    .B(_05086_),
    .X(_02684_));
 sky130_vsdinv _21720_ (.A(_05012_),
    .Y(_05087_));
 sky130_fd_sc_hd__o21ai_2 _21721_ (.A1(_05087_),
    .A2(_05079_),
    .B1(_05081_),
    .Y(_05088_));
 sky130_fd_sc_hd__clkbuf_4 _21722_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05089_));
 sky130_fd_sc_hd__clkbuf_4 _21723_ (.A(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__buf_4 _21724_ (.A(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__buf_6 _21725_ (.A(_05091_),
    .X(_05092_));
 sky130_fd_sc_hd__nor3_4 _21726_ (.A(_14086_),
    .B(_14435_),
    .C(_05043_),
    .Y(_05093_));
 sky130_fd_sc_hd__a41oi_4 _21727_ (.A1(_04946_),
    .A2(_04947_),
    .A3(_05092_),
    .A4(_05033_),
    .B1(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__nor2_1 _21728_ (.A(_05055_),
    .B(_05058_),
    .Y(_05095_));
 sky130_fd_sc_hd__o21bai_4 _21729_ (.A1(_05044_),
    .A2(_05059_),
    .B1_N(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__and2_2 _21730_ (.A(_14082_),
    .B(_05033_),
    .X(_05097_));
 sky130_fd_sc_hd__buf_4 _21731_ (.A(_14420_),
    .X(_05098_));
 sky130_fd_sc_hd__buf_4 _21732_ (.A(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__nand2_2 _21733_ (.A(_14090_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__clkbuf_4 _21734_ (.A(_05047_),
    .X(_05101_));
 sky130_fd_sc_hd__nand2_2 _21735_ (.A(_04909_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__xnor2_4 _21736_ (.A(_05100_),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__xor2_4 _21737_ (.A(_05097_),
    .B(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__buf_2 _21738_ (.A(_14408_),
    .X(_05105_));
 sky130_fd_sc_hd__buf_4 _21739_ (.A(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__nand2_2 _21740_ (.A(_05045_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__buf_4 _21741_ (.A(_04962_),
    .X(_05108_));
 sky130_fd_sc_hd__clkbuf_4 _21742_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05109_));
 sky130_fd_sc_hd__nand3_4 _21743_ (.A(_05108_),
    .B(_05109_),
    .C(_04956_),
    .Y(_05110_));
 sky130_fd_sc_hd__buf_4 _21744_ (.A(_04926_),
    .X(_05111_));
 sky130_fd_sc_hd__a22o_1 _21745_ (.A1(_14073_),
    .A2(_04897_),
    .B1(_05050_),
    .B2(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__o21ai_4 _21746_ (.A1(_14437_),
    .A2(_05110_),
    .B1(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__xnor2_4 _21747_ (.A(_05107_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__clkbuf_4 _21748_ (.A(_14416_),
    .X(_05115_));
 sky130_fd_sc_hd__clkbuf_4 _21749_ (.A(_04962_),
    .X(_05116_));
 sky130_fd_sc_hd__buf_4 _21750_ (.A(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__nand3b_1 _21751_ (.A_N(_05052_),
    .B(_05117_),
    .C(_04937_),
    .Y(_05118_));
 sky130_fd_sc_hd__o31a_2 _21752_ (.A1(_05056_),
    .A2(_05115_),
    .A3(_05054_),
    .B1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__xnor2_4 _21753_ (.A(_05114_),
    .B(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__xor2_4 _21754_ (.A(_05104_),
    .B(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__xnor2_2 _21755_ (.A(_05096_),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__xor2_2 _21756_ (.A(_05094_),
    .B(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__nor2_4 _21757_ (.A(_05066_),
    .B(_05067_),
    .Y(_05124_));
 sky130_fd_sc_hd__nand2_1 _21758_ (.A(_04999_),
    .B(_04891_),
    .Y(_05125_));
 sky130_fd_sc_hd__buf_6 _21759_ (.A(_14062_),
    .X(_05126_));
 sky130_fd_sc_hd__buf_6 _21760_ (.A(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__nand3_4 _21761_ (.A(_05127_),
    .B(_05065_),
    .C(_04908_),
    .Y(_05128_));
 sky130_fd_sc_hd__buf_2 _21762_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05129_));
 sky130_fd_sc_hd__clkbuf_4 _21763_ (.A(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__buf_6 _21764_ (.A(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__buf_4 _21765_ (.A(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__a22o_1 _21766_ (.A1(_05132_),
    .A2(_04717_),
    .B1(_05065_),
    .B2(_04872_),
    .X(_05133_));
 sky130_fd_sc_hd__o21ai_2 _21767_ (.A1(_14453_),
    .A2(_05128_),
    .B1(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__xnor2_1 _21768_ (.A(_05125_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__xnor2_1 _21769_ (.A(_05124_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__and2_1 _21770_ (.A(_05123_),
    .B(_05136_),
    .X(_05137_));
 sky130_vsdinv _21771_ (.A(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__or2_2 _21772_ (.A(_05136_),
    .B(_05123_),
    .X(_05139_));
 sky130_fd_sc_hd__a21o_1 _21773_ (.A1(_05138_),
    .A2(_05139_),
    .B1(_05070_),
    .X(_05140_));
 sky130_fd_sc_hd__nand3b_4 _21774_ (.A_N(_05137_),
    .B(_05070_),
    .C(_05139_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_1 _21775_ (.A(_05140_),
    .B(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__a21oi_4 _21776_ (.A1(_05060_),
    .A2(_05037_),
    .B1(_05062_),
    .Y(_05143_));
 sky130_fd_sc_hd__nor2_1 _21777_ (.A(_05143_),
    .B(_05075_),
    .Y(_05144_));
 sky130_vsdinv _21778_ (.A(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__nand2_1 _21779_ (.A(_05075_),
    .B(_05143_),
    .Y(_05146_));
 sky130_fd_sc_hd__nand3b_1 _21780_ (.A_N(_05142_),
    .B(_05145_),
    .C(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__xnor2_1 _21781_ (.A(_05143_),
    .B(_05075_),
    .Y(_05148_));
 sky130_fd_sc_hd__nand2_1 _21782_ (.A(_05148_),
    .B(_05142_),
    .Y(_05149_));
 sky130_fd_sc_hd__nand2_1 _21783_ (.A(_05147_),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__xnor2_2 _21784_ (.A(_05088_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__nor3b_1 _21785_ (.A(_05014_),
    .B(_05012_),
    .C_N(_05021_),
    .Y(_05152_));
 sky130_fd_sc_hd__nor3b_2 _21786_ (.A(_05079_),
    .B(_05082_),
    .C_N(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__a21o_1 _21787_ (.A1(_05086_),
    .A2(_05031_),
    .B1(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__xor2_1 _21788_ (.A(_05151_),
    .B(_05154_),
    .X(_02685_));
 sky130_fd_sc_hd__nor3b_1 _21789_ (.A(_05087_),
    .B(_05079_),
    .C_N(_05081_),
    .Y(_05155_));
 sky130_fd_sc_hd__and2b_1 _21790_ (.A_N(_05150_),
    .B(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__a21oi_4 _21791_ (.A1(_05154_),
    .A2(_05151_),
    .B1(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2b_4 _21792_ (.A_N(_05135_),
    .B(_05124_),
    .Y(_05158_));
 sky130_fd_sc_hd__o22a_2 _21793_ (.A1(_14454_),
    .A2(_05128_),
    .B1(_05125_),
    .B2(_05134_),
    .X(_05159_));
 sky130_fd_sc_hd__and2_2 _21794_ (.A(_04998_),
    .B(_04899_),
    .X(_05160_));
 sky130_fd_sc_hd__nand2_2 _21795_ (.A(_05126_),
    .B(_04907_),
    .Y(_05161_));
 sky130_fd_sc_hd__buf_6 _21796_ (.A(\pcpi_mul.rs2[7] ),
    .X(_05162_));
 sky130_fd_sc_hd__buf_6 _21797_ (.A(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__buf_6 _21798_ (.A(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__nand2_2 _21799_ (.A(_05164_),
    .B(_04969_),
    .Y(_05165_));
 sky130_fd_sc_hd__xnor2_4 _21800_ (.A(_05161_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__xor2_4 _21801_ (.A(_05160_),
    .B(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__xnor2_4 _21802_ (.A(_05159_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__xor2_1 _21803_ (.A(_05158_),
    .B(_05168_),
    .X(_05169_));
 sky130_vsdinv _21804_ (.A(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__nor2_1 _21805_ (.A(_05114_),
    .B(_05119_),
    .Y(_05171_));
 sky130_fd_sc_hd__o21bai_4 _21806_ (.A1(_05104_),
    .A2(_05120_),
    .B1_N(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__and2_2 _21807_ (.A(_14082_),
    .B(_05041_),
    .X(_05173_));
 sky130_fd_sc_hd__nand2_2 _21808_ (.A(_14090_),
    .B(_05048_),
    .Y(_05174_));
 sky130_fd_sc_hd__nand2_2 _21809_ (.A(_14093_),
    .B(_05106_),
    .Y(_05175_));
 sky130_fd_sc_hd__xnor2_4 _21810_ (.A(_05174_),
    .B(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__xor2_4 _21811_ (.A(_05173_),
    .B(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__buf_4 _21812_ (.A(_14438_),
    .X(_05178_));
 sky130_fd_sc_hd__o22a_2 _21813_ (.A1(_05178_),
    .A2(_05110_),
    .B1(_05107_),
    .B2(_05113_),
    .X(_05179_));
 sky130_fd_sc_hd__clkbuf_2 _21814_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_4 _21815_ (.A(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__and2_2 _21816_ (.A(_04712_),
    .B(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__nand2_2 _21817_ (.A(_04985_),
    .B(_14432_),
    .Y(_05183_));
 sky130_fd_sc_hd__clkbuf_4 _21818_ (.A(_04959_),
    .X(_05184_));
 sky130_fd_sc_hd__nand2_2 _21819_ (.A(_04923_),
    .B(_05184_),
    .Y(_05185_));
 sky130_fd_sc_hd__xnor2_4 _21820_ (.A(_05183_),
    .B(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__xor2_4 _21821_ (.A(_05182_),
    .B(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__xnor2_4 _21822_ (.A(_05179_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__xor2_4 _21823_ (.A(_05177_),
    .B(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__xor2_1 _21824_ (.A(_05172_),
    .B(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__buf_4 _21825_ (.A(_05101_),
    .X(_05191_));
 sky130_fd_sc_hd__nor3_4 _21826_ (.A(_14085_),
    .B(_14429_),
    .C(_05103_),
    .Y(_05192_));
 sky130_fd_sc_hd__a41oi_4 _21827_ (.A1(_04886_),
    .A2(_04878_),
    .A3(_05191_),
    .A4(_05092_),
    .B1(_05192_),
    .Y(_05193_));
 sky130_vsdinv _21828_ (.A(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__and2_2 _21829_ (.A(_05190_),
    .B(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__or2b_1 _21830_ (.A(_05190_),
    .B_N(_05193_),
    .X(_05196_));
 sky130_fd_sc_hd__nor3b_4 _21831_ (.A(_05170_),
    .B(_05195_),
    .C_N(_05196_),
    .Y(_05197_));
 sky130_vsdinv _21832_ (.A(_05197_),
    .Y(_05198_));
 sky130_vsdinv _21833_ (.A(_05195_),
    .Y(_05199_));
 sky130_fd_sc_hd__a21o_1 _21834_ (.A1(_05199_),
    .A2(_05196_),
    .B1(_05169_),
    .X(_05200_));
 sky130_fd_sc_hd__and3_4 _21835_ (.A(_05137_),
    .B(_05198_),
    .C(_05200_),
    .X(_05201_));
 sky130_vsdinv _21836_ (.A(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__a21o_1 _21837_ (.A1(_05198_),
    .A2(_05200_),
    .B1(_05137_),
    .X(_05203_));
 sky130_fd_sc_hd__buf_2 _21838_ (.A(\pcpi_mul.rs2[9] ),
    .X(_05204_));
 sky130_fd_sc_hd__buf_2 _21839_ (.A(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__buf_4 _21840_ (.A(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__and2_1 _21841_ (.A(_05206_),
    .B(_04721_),
    .X(_05207_));
 sky130_fd_sc_hd__a21oi_2 _21842_ (.A1(_05202_),
    .A2(_05203_),
    .B1(_05207_),
    .Y(_05208_));
 sky130_vsdinv _21843_ (.A(_05207_),
    .Y(_05209_));
 sky130_fd_sc_hd__nor3b_4 _21844_ (.A(_05209_),
    .B(_05201_),
    .C_N(_05203_),
    .Y(_05210_));
 sky130_vsdinv _21845_ (.A(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__nor2_2 _21846_ (.A(_05094_),
    .B(_05122_),
    .Y(_05212_));
 sky130_fd_sc_hd__a21oi_4 _21847_ (.A1(_05121_),
    .A2(_05096_),
    .B1(_05212_),
    .Y(_05213_));
 sky130_fd_sc_hd__xor2_4 _21848_ (.A(_05213_),
    .B(_05141_),
    .X(_05214_));
 sky130_fd_sc_hd__nand3b_4 _21849_ (.A_N(_05208_),
    .B(_05211_),
    .C(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__o21bai_2 _21850_ (.A1(_05210_),
    .A2(_05208_),
    .B1_N(_05214_),
    .Y(_05216_));
 sky130_fd_sc_hd__a31oi_1 _21851_ (.A1(_05140_),
    .A2(_05146_),
    .A3(_05141_),
    .B1(_05144_),
    .Y(_05217_));
 sky130_vsdinv _21852_ (.A(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__a21oi_2 _21853_ (.A1(_05215_),
    .A2(_05216_),
    .B1(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__nand3_4 _21854_ (.A(_05215_),
    .B(_05216_),
    .C(_05218_),
    .Y(_05220_));
 sky130_vsdinv _21855_ (.A(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__and3_1 _21856_ (.A(_05147_),
    .B(_05149_),
    .C(_05082_),
    .X(_05222_));
 sky130_fd_sc_hd__nor3b_2 _21857_ (.A(_05219_),
    .B(_05221_),
    .C_N(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__o21ba_1 _21858_ (.A1(_05219_),
    .A2(_05221_),
    .B1_N(_05222_),
    .X(_05224_));
 sky130_fd_sc_hd__nor2_1 _21859_ (.A(_05223_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__xnor2_1 _21860_ (.A(_05157_),
    .B(_05225_),
    .Y(_02686_));
 sky130_fd_sc_hd__o21bai_2 _21861_ (.A1(_05224_),
    .A2(_05157_),
    .B1_N(_05223_),
    .Y(_05226_));
 sky130_fd_sc_hd__buf_4 _21862_ (.A(_14408_),
    .X(_05227_));
 sky130_fd_sc_hd__buf_4 _21863_ (.A(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__buf_4 _21864_ (.A(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__nor3_4 _21865_ (.A(_14086_),
    .B(_14423_),
    .C(_05176_),
    .Y(_05230_));
 sky130_fd_sc_hd__a41oi_4 _21866_ (.A1(_04946_),
    .A2(_04879_),
    .A3(_05229_),
    .A4(_05191_),
    .B1(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__nor2_1 _21867_ (.A(_05179_),
    .B(_05187_),
    .Y(_05232_));
 sky130_fd_sc_hd__o21bai_4 _21868_ (.A1(_05177_),
    .A2(_05188_),
    .B1_N(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__and2_2 _21869_ (.A(_04932_),
    .B(_05191_),
    .X(_05234_));
 sky130_fd_sc_hd__nand2_2 _21870_ (.A(_04904_),
    .B(_05228_),
    .Y(_05235_));
 sky130_fd_sc_hd__buf_2 _21871_ (.A(_05180_),
    .X(_05236_));
 sky130_fd_sc_hd__buf_4 _21872_ (.A(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__nand2_2 _21873_ (.A(_04909_),
    .B(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__xnor2_4 _21874_ (.A(_05235_),
    .B(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__xor2_4 _21875_ (.A(_05234_),
    .B(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__buf_2 _21876_ (.A(_14398_),
    .X(_05241_));
 sky130_fd_sc_hd__and2_2 _21877_ (.A(_05045_),
    .B(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__nand2_2 _21878_ (.A(_05109_),
    .B(_05098_),
    .Y(_05243_));
 sky130_fd_sc_hd__and2_1 _21879_ (.A(_04962_),
    .B(_05184_),
    .X(_05244_));
 sky130_fd_sc_hd__xor2_4 _21880_ (.A(_05243_),
    .B(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__xor2_4 _21881_ (.A(_05242_),
    .B(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__buf_6 _21882_ (.A(_14428_),
    .X(_05247_));
 sky130_fd_sc_hd__o32a_4 _21883_ (.A1(_05056_),
    .A2(_14405_),
    .A3(_05186_),
    .B1(_05247_),
    .B2(_05110_),
    .X(_05248_));
 sky130_fd_sc_hd__xnor2_4 _21884_ (.A(_05246_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__xor2_4 _21885_ (.A(_05240_),
    .B(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__xnor2_2 _21886_ (.A(_05233_),
    .B(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__nor2_4 _21887_ (.A(_05231_),
    .B(_05251_),
    .Y(_05252_));
 sky130_vsdinv _21888_ (.A(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2_1 _21889_ (.A(_05251_),
    .B(_05231_),
    .Y(_05254_));
 sky130_fd_sc_hd__and2_2 _21890_ (.A(_04999_),
    .B(_04929_),
    .X(_05255_));
 sky130_fd_sc_hd__nand2_2 _21891_ (.A(_05065_),
    .B(_04899_),
    .Y(_05256_));
 sky130_fd_sc_hd__and2_1 _21892_ (.A(_05132_),
    .B(_04969_),
    .X(_05257_));
 sky130_fd_sc_hd__xor2_4 _21893_ (.A(_05256_),
    .B(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__xor2_4 _21894_ (.A(_05255_),
    .B(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__o32a_4 _21895_ (.A1(_14071_),
    .A2(_14439_),
    .A3(_05166_),
    .B1(_14445_),
    .B2(_05128_),
    .X(_05260_));
 sky130_fd_sc_hd__xnor2_4 _21896_ (.A(_05259_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__or2_4 _21897_ (.A(_05159_),
    .B(_05167_),
    .X(_05262_));
 sky130_fd_sc_hd__o21ai_4 _21898_ (.A1(_05158_),
    .A2(_05168_),
    .B1(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__xor2_4 _21899_ (.A(_05261_),
    .B(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__a21boi_2 _21900_ (.A1(_05253_),
    .A2(_05254_),
    .B1_N(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__nor3b_4 _21901_ (.A(_05264_),
    .B(_05252_),
    .C_N(_05254_),
    .Y(_05266_));
 sky130_vsdinv _21902_ (.A(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand3b_4 _21903_ (.A_N(_05265_),
    .B(_05197_),
    .C(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__o21bai_2 _21904_ (.A1(_05266_),
    .A2(_05265_),
    .B1_N(_05197_),
    .Y(_05269_));
 sky130_fd_sc_hd__or4_4 _21905_ (.A(_14054_),
    .B(_14059_),
    .C(_14449_),
    .D(_14453_),
    .X(_05270_));
 sky130_fd_sc_hd__buf_6 _21906_ (.A(\pcpi_mul.rs2[10] ),
    .X(_05271_));
 sky130_fd_sc_hd__clkbuf_4 _21907_ (.A(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__buf_6 _21908_ (.A(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__buf_6 _21909_ (.A(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__a22o_1 _21910_ (.A1(_05274_),
    .A2(_04721_),
    .B1(_05206_),
    .B2(_04874_),
    .X(_05275_));
 sky130_fd_sc_hd__and2_1 _21911_ (.A(_05270_),
    .B(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__and3_2 _21912_ (.A(_05268_),
    .B(_05269_),
    .C(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__a21oi_4 _21913_ (.A1(_05268_),
    .A2(_05269_),
    .B1(_05276_),
    .Y(_05278_));
 sky130_fd_sc_hd__nor3b_4 _21914_ (.A(_05277_),
    .B(_05278_),
    .C_N(_05210_),
    .Y(_05279_));
 sky130_vsdinv _21915_ (.A(_05277_),
    .Y(_05280_));
 sky130_vsdinv _21916_ (.A(_05278_),
    .Y(_05281_));
 sky130_fd_sc_hd__a21oi_2 _21917_ (.A1(_05280_),
    .A2(_05281_),
    .B1(_05210_),
    .Y(_05282_));
 sky130_vsdinv _21918_ (.A(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__a21oi_4 _21919_ (.A1(_05189_),
    .A2(_05172_),
    .B1(_05195_),
    .Y(_05284_));
 sky130_vsdinv _21920_ (.A(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__xor2_4 _21921_ (.A(_05285_),
    .B(_05201_),
    .X(_05286_));
 sky130_fd_sc_hd__nand3b_4 _21922_ (.A_N(_05279_),
    .B(_05283_),
    .C(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__o21bai_2 _21923_ (.A1(_05282_),
    .A2(_05279_),
    .B1_N(_05286_),
    .Y(_05288_));
 sky130_fd_sc_hd__o21a_2 _21924_ (.A1(_05141_),
    .A2(_05213_),
    .B1(_05215_),
    .X(_05289_));
 sky130_fd_sc_hd__a21boi_4 _21925_ (.A1(_05287_),
    .A2(_05288_),
    .B1_N(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand2_2 _21926_ (.A(_05287_),
    .B(_05288_),
    .Y(_05291_));
 sky130_fd_sc_hd__nor2_8 _21927_ (.A(_05289_),
    .B(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__nor3_4 _21928_ (.A(_05220_),
    .B(_05290_),
    .C(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__o21bai_2 _21929_ (.A1(_05290_),
    .A2(_05292_),
    .B1_N(_05221_),
    .Y(_05294_));
 sky130_fd_sc_hd__and2b_1 _21930_ (.A_N(_05293_),
    .B(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__xor2_1 _21931_ (.A(_05226_),
    .B(_05295_),
    .X(_02629_));
 sky130_fd_sc_hd__a21oi_4 _21932_ (.A1(_05226_),
    .A2(_05294_),
    .B1(_05293_),
    .Y(_05296_));
 sky130_fd_sc_hd__a21o_1 _21933_ (.A1(_05283_),
    .A2(_05286_),
    .B1(_05279_),
    .X(_05297_));
 sky130_fd_sc_hd__buf_6 _21934_ (.A(_04886_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_8 _21935_ (.A(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__buf_6 _21936_ (.A(_04947_),
    .X(_05300_));
 sky130_fd_sc_hd__buf_4 _21937_ (.A(_05237_),
    .X(_05301_));
 sky130_fd_sc_hd__clkbuf_8 _21938_ (.A(_14086_),
    .X(_05302_));
 sky130_fd_sc_hd__nor3_4 _21939_ (.A(_05302_),
    .B(_14418_),
    .C(_05239_),
    .Y(_05303_));
 sky130_fd_sc_hd__a41oi_4 _21940_ (.A1(_05299_),
    .A2(_05300_),
    .A3(_05301_),
    .A4(_05229_),
    .B1(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__nor2_1 _21941_ (.A(_05246_),
    .B(_05248_),
    .Y(_05305_));
 sky130_fd_sc_hd__o21bai_4 _21942_ (.A1(_05240_),
    .A2(_05249_),
    .B1_N(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__and2_2 _21943_ (.A(_04933_),
    .B(_05229_),
    .X(_05307_));
 sky130_fd_sc_hd__clkbuf_4 _21944_ (.A(_05180_),
    .X(_05308_));
 sky130_fd_sc_hd__buf_4 _21945_ (.A(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__nand2_2 _21946_ (.A(_04905_),
    .B(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__buf_4 _21947_ (.A(_05241_),
    .X(_05311_));
 sky130_fd_sc_hd__nand2_2 _21948_ (.A(_04910_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__xnor2_4 _21949_ (.A(_05310_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__xor2_4 _21950_ (.A(_05307_),
    .B(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__clkbuf_4 _21951_ (.A(_14096_),
    .X(_05315_));
 sky130_fd_sc_hd__buf_4 _21952_ (.A(_05117_),
    .X(_05316_));
 sky130_fd_sc_hd__nand3b_1 _21953_ (.A_N(_05243_),
    .B(_05316_),
    .C(_05033_),
    .Y(_05317_));
 sky130_fd_sc_hd__o31a_2 _21954_ (.A1(_05315_),
    .A2(_14401_),
    .A3(_05245_),
    .B1(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__buf_4 _21955_ (.A(_04712_),
    .X(_05319_));
 sky130_fd_sc_hd__clkbuf_2 _21956_ (.A(\pcpi_mul.rs1[11] ),
    .X(_05320_));
 sky130_fd_sc_hd__buf_2 _21957_ (.A(_05320_),
    .X(_05321_));
 sky130_fd_sc_hd__clkbuf_4 _21958_ (.A(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__and2_2 _21959_ (.A(_05319_),
    .B(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__buf_6 _21960_ (.A(_05050_),
    .X(_05324_));
 sky130_fd_sc_hd__nand2_2 _21961_ (.A(_05324_),
    .B(_05048_),
    .Y(_05325_));
 sky130_fd_sc_hd__clkbuf_4 _21962_ (.A(_04962_),
    .X(_05326_));
 sky130_fd_sc_hd__and2_1 _21963_ (.A(_05326_),
    .B(_04983_),
    .X(_05327_));
 sky130_fd_sc_hd__xor2_4 _21964_ (.A(_05325_),
    .B(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__xor2_4 _21965_ (.A(_05323_),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__xnor2_4 _21966_ (.A(_05318_),
    .B(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__xor2_4 _21967_ (.A(_05314_),
    .B(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__xnor2_2 _21968_ (.A(_05306_),
    .B(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__nor2_2 _21969_ (.A(_05304_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__nand2_2 _21970_ (.A(_05332_),
    .B(_05304_),
    .Y(_05334_));
 sky130_fd_sc_hd__nor2_2 _21971_ (.A(_05259_),
    .B(_05260_),
    .Y(_05335_));
 sky130_fd_sc_hd__o21bai_4 _21972_ (.A1(_05262_),
    .A2(_05261_),
    .B1_N(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__buf_6 _21973_ (.A(_05127_),
    .X(_05337_));
 sky130_fd_sc_hd__nand3b_2 _21974_ (.A_N(_05256_),
    .B(_05337_),
    .C(_04891_),
    .Y(_05338_));
 sky130_fd_sc_hd__o31a_4 _21975_ (.A1(_14071_),
    .A2(_14435_),
    .A3(_05258_),
    .B1(_05338_),
    .X(_05339_));
 sky130_fd_sc_hd__and2_2 _21976_ (.A(_04998_),
    .B(_05039_),
    .X(_05340_));
 sky130_fd_sc_hd__nand2_2 _21977_ (.A(_05164_),
    .B(_04976_),
    .Y(_05341_));
 sky130_fd_sc_hd__and2_1 _21978_ (.A(_05131_),
    .B(_04949_),
    .X(_05342_));
 sky130_fd_sc_hd__xor2_4 _21979_ (.A(_05341_),
    .B(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__xor2_4 _21980_ (.A(_05340_),
    .B(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__xnor2_4 _21981_ (.A(_05270_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__xor2_4 _21982_ (.A(_05339_),
    .B(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__xor2_4 _21983_ (.A(_05336_),
    .B(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__nand3b_4 _21984_ (.A_N(_05333_),
    .B(_05334_),
    .C(_05347_),
    .Y(_05348_));
 sky130_vsdinv _21985_ (.A(_05333_),
    .Y(_05349_));
 sky130_fd_sc_hd__a21o_1 _21986_ (.A1(_05349_),
    .A2(_05334_),
    .B1(_05347_),
    .X(_05350_));
 sky130_fd_sc_hd__o31ai_4 _21987_ (.A1(_05158_),
    .A2(_05168_),
    .A3(_05261_),
    .B1(_05267_),
    .Y(_05351_));
 sky130_fd_sc_hd__a21o_1 _21988_ (.A1(_05348_),
    .A2(_05350_),
    .B1(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__nand3_4 _21989_ (.A(_05351_),
    .B(_05350_),
    .C(_05348_),
    .Y(_05353_));
 sky130_fd_sc_hd__buf_2 _21990_ (.A(\pcpi_mul.rs2[9] ),
    .X(_05354_));
 sky130_fd_sc_hd__clkbuf_4 _21991_ (.A(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__and2_2 _21992_ (.A(_05355_),
    .B(_04937_),
    .X(_05356_));
 sky130_fd_sc_hd__buf_2 _21993_ (.A(\pcpi_mul.rs2[11] ),
    .X(_05357_));
 sky130_fd_sc_hd__buf_4 _21994_ (.A(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__buf_6 _21995_ (.A(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__nand3_4 _21996_ (.A(_05359_),
    .B(_05273_),
    .C(_04907_),
    .Y(_05360_));
 sky130_fd_sc_hd__buf_4 _21997_ (.A(_14050_),
    .X(_05361_));
 sky130_fd_sc_hd__buf_4 _21998_ (.A(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__buf_4 _21999_ (.A(_05272_),
    .X(_05363_));
 sky130_fd_sc_hd__buf_4 _22000_ (.A(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__a22o_2 _22001_ (.A1(_05362_),
    .A2(_04717_),
    .B1(_05364_),
    .B2(_04908_),
    .X(_05365_));
 sky130_fd_sc_hd__o21ai_4 _22002_ (.A1(_14454_),
    .A2(_05360_),
    .B1(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__xnor2_4 _22003_ (.A(_05356_),
    .B(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__a21o_1 _22004_ (.A1(_05352_),
    .A2(_05353_),
    .B1(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__nand3_4 _22005_ (.A(_05352_),
    .B(_05367_),
    .C(_05353_),
    .Y(_05369_));
 sky130_fd_sc_hd__a21oi_2 _22006_ (.A1(_05368_),
    .A2(_05369_),
    .B1(_05277_),
    .Y(_05370_));
 sky130_fd_sc_hd__a21oi_4 _22007_ (.A1(_05250_),
    .A2(_05233_),
    .B1(_05252_),
    .Y(_05371_));
 sky130_fd_sc_hd__xor2_4 _22008_ (.A(_05371_),
    .B(_05268_),
    .X(_05372_));
 sky130_fd_sc_hd__nand3_4 _22009_ (.A(_05368_),
    .B(_05277_),
    .C(_05369_),
    .Y(_05373_));
 sky130_fd_sc_hd__nand3b_4 _22010_ (.A_N(_05370_),
    .B(_05372_),
    .C(_05373_),
    .Y(_05374_));
 sky130_vsdinv _22011_ (.A(_05373_),
    .Y(_05375_));
 sky130_fd_sc_hd__o21bai_2 _22012_ (.A1(_05370_),
    .A2(_05375_),
    .B1_N(_05372_),
    .Y(_05376_));
 sky130_fd_sc_hd__nand3_4 _22013_ (.A(_05297_),
    .B(_05374_),
    .C(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__a21o_1 _22014_ (.A1(_05376_),
    .A2(_05374_),
    .B1(_05297_),
    .X(_05378_));
 sky130_fd_sc_hd__o2bb2ai_1 _22015_ (.A1_N(_05377_),
    .A2_N(_05378_),
    .B1(_05202_),
    .B2(_05284_),
    .Y(_05379_));
 sky130_fd_sc_hd__and4_2 _22016_ (.A(_05137_),
    .B(_05198_),
    .C(_05200_),
    .D(_05285_),
    .X(_05380_));
 sky130_fd_sc_hd__nand3_2 _22017_ (.A(_05378_),
    .B(_05380_),
    .C(_05377_),
    .Y(_05381_));
 sky130_fd_sc_hd__a21oi_2 _22018_ (.A1(_05379_),
    .A2(_05381_),
    .B1(_05292_),
    .Y(_05382_));
 sky130_vsdinv _22019_ (.A(_05292_),
    .Y(_05383_));
 sky130_fd_sc_hd__a21oi_1 _22020_ (.A1(_05378_),
    .A2(_05377_),
    .B1(_05380_),
    .Y(_05384_));
 sky130_fd_sc_hd__nor3b_2 _22021_ (.A(_05383_),
    .B(_05384_),
    .C_N(_05381_),
    .Y(_05385_));
 sky130_fd_sc_hd__nor2_1 _22022_ (.A(_05382_),
    .B(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__xnor2_1 _22023_ (.A(_05296_),
    .B(_05386_),
    .Y(_02630_));
 sky130_fd_sc_hd__or3b_4 _22024_ (.A(_05262_),
    .B(_05261_),
    .C_N(_05346_),
    .X(_05387_));
 sky130_fd_sc_hd__nand2_4 _22025_ (.A(_05346_),
    .B(_05335_),
    .Y(_05388_));
 sky130_fd_sc_hd__or2_1 _22026_ (.A(_05270_),
    .B(_05344_),
    .X(_05389_));
 sky130_fd_sc_hd__o21ai_4 _22027_ (.A1(_05339_),
    .A2(_05345_),
    .B1(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__nand3b_1 _22028_ (.A_N(_05341_),
    .B(_05337_),
    .C(_04900_),
    .Y(_05391_));
 sky130_fd_sc_hd__o31a_2 _22029_ (.A1(_14071_),
    .A2(_14429_),
    .A3(_05343_),
    .B1(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__a2bb2oi_4 _22030_ (.A1_N(_14454_),
    .A2_N(_05360_),
    .B1(_05356_),
    .B2(_05365_),
    .Y(_05393_));
 sky130_fd_sc_hd__and2_2 _22031_ (.A(_04997_),
    .B(_05041_),
    .X(_05394_));
 sky130_fd_sc_hd__nand2_2 _22032_ (.A(_05064_),
    .B(_04978_),
    .Y(_05395_));
 sky130_fd_sc_hd__and2_1 _22033_ (.A(_05131_),
    .B(_04927_),
    .X(_05396_));
 sky130_fd_sc_hd__xor2_4 _22034_ (.A(_05395_),
    .B(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__xor2_4 _22035_ (.A(_05394_),
    .B(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__xnor2_4 _22036_ (.A(_05393_),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__xor2_4 _22037_ (.A(_05392_),
    .B(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__xnor2_4 _22038_ (.A(_05390_),
    .B(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__xor2_4 _22039_ (.A(_05388_),
    .B(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__buf_6 _22040_ (.A(_04946_),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_4 _22041_ (.A(_14398_),
    .X(_05404_));
 sky130_fd_sc_hd__buf_4 _22042_ (.A(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__buf_4 _22043_ (.A(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__nor3_4 _22044_ (.A(_14087_),
    .B(_14412_),
    .C(_05313_),
    .Y(_05407_));
 sky130_fd_sc_hd__a41oi_4 _22045_ (.A1(_05403_),
    .A2(_05300_),
    .A3(_05406_),
    .A4(_05301_),
    .B1(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__nor2_1 _22046_ (.A(_05318_),
    .B(_05329_),
    .Y(_05409_));
 sky130_fd_sc_hd__o21bai_4 _22047_ (.A1(_05314_),
    .A2(_05330_),
    .B1_N(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__and2_2 _22048_ (.A(_14083_),
    .B(_05301_),
    .X(_05411_));
 sky130_fd_sc_hd__nand2_2 _22049_ (.A(_04936_),
    .B(_05311_),
    .Y(_05412_));
 sky130_fd_sc_hd__buf_2 _22050_ (.A(_05320_),
    .X(_05413_));
 sky130_fd_sc_hd__buf_4 _22051_ (.A(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__nand2_2 _22052_ (.A(_04910_),
    .B(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__xnor2_4 _22053_ (.A(_05412_),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__xor2_4 _22054_ (.A(_05411_),
    .B(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__buf_6 _22055_ (.A(_14394_),
    .X(_05418_));
 sky130_fd_sc_hd__clkbuf_4 _22056_ (.A(_04985_),
    .X(_05419_));
 sky130_fd_sc_hd__clkbuf_4 _22057_ (.A(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__nand3b_1 _22058_ (.A_N(_05325_),
    .B(_05420_),
    .C(_05092_),
    .Y(_05421_));
 sky130_fd_sc_hd__o31a_2 _22059_ (.A1(_05315_),
    .A2(_05418_),
    .A3(_05328_),
    .B1(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__clkbuf_4 _22060_ (.A(_14387_),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_4 _22061_ (.A(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__and2_2 _22062_ (.A(_04955_),
    .B(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_2 _22063_ (.A(_14408_),
    .X(_05426_));
 sky130_fd_sc_hd__clkbuf_4 _22064_ (.A(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__nand2_2 _22065_ (.A(_05324_),
    .B(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__buf_4 _22066_ (.A(_05046_),
    .X(_05429_));
 sky130_fd_sc_hd__and2_1 _22067_ (.A(_05326_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__xor2_4 _22068_ (.A(_05428_),
    .B(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__xor2_4 _22069_ (.A(_05425_),
    .B(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__xnor2_4 _22070_ (.A(_05422_),
    .B(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__xor2_4 _22071_ (.A(_05417_),
    .B(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__xnor2_4 _22072_ (.A(_05410_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__xor2_4 _22073_ (.A(_05408_),
    .B(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__xnor2_4 _22074_ (.A(_05402_),
    .B(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__a21o_2 _22075_ (.A1(_05348_),
    .A2(_05387_),
    .B1(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__nand3_4 _22076_ (.A(_05437_),
    .B(_05348_),
    .C(_05387_),
    .Y(_05439_));
 sky130_fd_sc_hd__clkbuf_4 _22077_ (.A(\pcpi_mul.rs2[12] ),
    .X(_05440_));
 sky130_fd_sc_hd__buf_4 _22078_ (.A(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__buf_8 _22079_ (.A(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__and2_2 _22080_ (.A(_05442_),
    .B(_04721_),
    .X(_05443_));
 sky130_fd_sc_hd__and2_2 _22081_ (.A(_05355_),
    .B(_04899_),
    .X(_05444_));
 sky130_fd_sc_hd__buf_6 _22082_ (.A(_05357_),
    .X(_05445_));
 sky130_fd_sc_hd__nand2_2 _22083_ (.A(_05445_),
    .B(_04906_),
    .Y(_05446_));
 sky130_fd_sc_hd__clkbuf_4 _22084_ (.A(_05271_),
    .X(_05447_));
 sky130_fd_sc_hd__nand2_2 _22085_ (.A(_05447_),
    .B(_04889_),
    .Y(_05448_));
 sky130_fd_sc_hd__xnor2_4 _22086_ (.A(_05446_),
    .B(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__xor2_4 _22087_ (.A(_05444_),
    .B(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__xnor2_4 _22088_ (.A(_05443_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__a21o_1 _22089_ (.A1(_05438_),
    .A2(_05439_),
    .B1(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__nand3_4 _22090_ (.A(_05438_),
    .B(_05451_),
    .C(_05439_),
    .Y(_05453_));
 sky130_vsdinv _22091_ (.A(_05369_),
    .Y(_05454_));
 sky130_fd_sc_hd__a21oi_2 _22092_ (.A1(_05452_),
    .A2(_05453_),
    .B1(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand3_4 _22093_ (.A(_05452_),
    .B(_05454_),
    .C(_05453_),
    .Y(_05456_));
 sky130_vsdinv _22094_ (.A(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__a21o_1 _22095_ (.A1(_05331_),
    .A2(_05306_),
    .B1(_05333_),
    .X(_05458_));
 sky130_fd_sc_hd__xnor2_2 _22096_ (.A(_05458_),
    .B(_05353_),
    .Y(_05459_));
 sky130_fd_sc_hd__o21bai_2 _22097_ (.A1(_05455_),
    .A2(_05457_),
    .B1_N(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__nand3b_4 _22098_ (.A_N(_05455_),
    .B(_05456_),
    .C(_05459_),
    .Y(_05461_));
 sky130_fd_sc_hd__nand2_2 _22099_ (.A(_05374_),
    .B(_05373_),
    .Y(_05462_));
 sky130_fd_sc_hd__a21oi_1 _22100_ (.A1(_05460_),
    .A2(_05461_),
    .B1(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__nand3_4 _22101_ (.A(_05462_),
    .B(_05460_),
    .C(_05461_),
    .Y(_05464_));
 sky130_vsdinv _22102_ (.A(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__nor2_4 _22103_ (.A(_05371_),
    .B(_05268_),
    .Y(_05466_));
 sky130_fd_sc_hd__o21bai_1 _22104_ (.A1(_05463_),
    .A2(_05465_),
    .B1_N(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__a21o_1 _22105_ (.A1(_05460_),
    .A2(_05461_),
    .B1(_05462_),
    .X(_05468_));
 sky130_fd_sc_hd__nand3_2 _22106_ (.A(_05468_),
    .B(_05466_),
    .C(_05464_),
    .Y(_05469_));
 sky130_fd_sc_hd__a21boi_4 _22107_ (.A1(_05378_),
    .A2(_05380_),
    .B1_N(_05377_),
    .Y(_05470_));
 sky130_fd_sc_hd__a21boi_2 _22108_ (.A1(_05467_),
    .A2(_05469_),
    .B1_N(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__a21oi_2 _22109_ (.A1(_05468_),
    .A2(_05464_),
    .B1(_05466_),
    .Y(_05472_));
 sky130_fd_sc_hd__nor3b_4 _22110_ (.A(_05470_),
    .B(_05472_),
    .C_N(_05469_),
    .Y(_05473_));
 sky130_fd_sc_hd__nor2_4 _22111_ (.A(_05471_),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__o21bai_2 _22112_ (.A1(_05382_),
    .A2(_05296_),
    .B1_N(_05385_),
    .Y(_05475_));
 sky130_fd_sc_hd__xor2_1 _22113_ (.A(_05474_),
    .B(_05475_),
    .X(_02631_));
 sky130_fd_sc_hd__nor2_2 _22114_ (.A(_05388_),
    .B(_05401_),
    .Y(_05476_));
 sky130_fd_sc_hd__a21oi_4 _22115_ (.A1(_05436_),
    .A2(_05402_),
    .B1(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__nor2_1 _22116_ (.A(_05393_),
    .B(_05398_),
    .Y(_05478_));
 sky130_fd_sc_hd__o21ba_1 _22117_ (.A1(_05392_),
    .A2(_05399_),
    .B1_N(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__nand3b_4 _22118_ (.A_N(_05450_),
    .B(_05442_),
    .C(_04719_),
    .Y(_05480_));
 sky130_fd_sc_hd__nand3b_1 _22119_ (.A_N(_05395_),
    .B(_05337_),
    .C(_04929_),
    .Y(_05481_));
 sky130_fd_sc_hd__o31a_2 _22120_ (.A1(_14071_),
    .A2(_14423_),
    .A3(_05397_),
    .B1(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_4 _22121_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05483_));
 sky130_fd_sc_hd__and2_2 _22122_ (.A(_05483_),
    .B(_05048_),
    .X(_05484_));
 sky130_fd_sc_hd__nand2_2 _22123_ (.A(_05163_),
    .B(_05098_),
    .Y(_05485_));
 sky130_fd_sc_hd__clkbuf_4 _22124_ (.A(_05129_),
    .X(_05486_));
 sky130_fd_sc_hd__and2_1 _22125_ (.A(_05486_),
    .B(_05184_),
    .X(_05487_));
 sky130_fd_sc_hd__xor2_4 _22126_ (.A(_05485_),
    .B(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__xor2_4 _22127_ (.A(_05484_),
    .B(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__o32a_4 _22128_ (.A1(_14059_),
    .A2(_05178_),
    .A3(_05449_),
    .B1(_14444_),
    .B2(_05360_),
    .X(_05490_));
 sky130_fd_sc_hd__xnor2_4 _22129_ (.A(_05489_),
    .B(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__xor2_4 _22130_ (.A(_05482_),
    .B(_05491_),
    .X(_05492_));
 sky130_fd_sc_hd__xor2_4 _22131_ (.A(_05480_),
    .B(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__xor2_2 _22132_ (.A(_05479_),
    .B(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__a21o_1 _22133_ (.A1(_05400_),
    .A2(_05390_),
    .B1(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__nand3_2 _22134_ (.A(_05494_),
    .B(_05400_),
    .C(_05390_),
    .Y(_05496_));
 sky130_fd_sc_hd__clkbuf_4 _22135_ (.A(_05321_),
    .X(_05497_));
 sky130_fd_sc_hd__buf_4 _22136_ (.A(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__nor3_4 _22137_ (.A(_14087_),
    .B(_14406_),
    .C(_05416_),
    .Y(_05499_));
 sky130_fd_sc_hd__a41oi_4 _22138_ (.A1(_05403_),
    .A2(_05300_),
    .A3(_05498_),
    .A4(_05406_),
    .B1(_05499_),
    .Y(_05500_));
 sky130_fd_sc_hd__nor2_1 _22139_ (.A(_05422_),
    .B(_05432_),
    .Y(_05501_));
 sky130_fd_sc_hd__o21bai_4 _22140_ (.A1(_05417_),
    .A2(_05433_),
    .B1_N(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__and2_2 _22141_ (.A(_04933_),
    .B(_05406_),
    .X(_05503_));
 sky130_fd_sc_hd__nand2_2 _22142_ (.A(_04905_),
    .B(_05498_),
    .Y(_05504_));
 sky130_fd_sc_hd__buf_4 _22143_ (.A(_05423_),
    .X(_05505_));
 sky130_fd_sc_hd__nand2_2 _22144_ (.A(_04910_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__xnor2_4 _22145_ (.A(_05504_),
    .B(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__xor2_4 _22146_ (.A(_05503_),
    .B(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__nand3b_1 _22147_ (.A_N(_05428_),
    .B(_05420_),
    .C(_05191_),
    .Y(_05509_));
 sky130_fd_sc_hd__o31a_2 _22148_ (.A1(_05315_),
    .A2(_14390_),
    .A3(_05431_),
    .B1(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__clkbuf_4 _22149_ (.A(\pcpi_mul.rs1[13] ),
    .X(_05511_));
 sky130_fd_sc_hd__buf_4 _22150_ (.A(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__buf_2 _22151_ (.A(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__and2_2 _22152_ (.A(_05319_),
    .B(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__buf_4 _22153_ (.A(_05109_),
    .X(_05515_));
 sky130_fd_sc_hd__buf_4 _22154_ (.A(_05236_),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_2 _22155_ (.A(_05515_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__and2_1 _22156_ (.A(_05116_),
    .B(_05427_),
    .X(_05518_));
 sky130_fd_sc_hd__xor2_4 _22157_ (.A(_05517_),
    .B(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__xor2_4 _22158_ (.A(_05514_),
    .B(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__xnor2_4 _22159_ (.A(_05510_),
    .B(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__xor2_4 _22160_ (.A(_05508_),
    .B(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__xnor2_4 _22161_ (.A(_05502_),
    .B(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__xor2_4 _22162_ (.A(_05500_),
    .B(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__a21o_1 _22163_ (.A1(_05495_),
    .A2(_05496_),
    .B1(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__nand3_2 _22164_ (.A(_05495_),
    .B(_05524_),
    .C(_05496_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_4 _22165_ (.A(_05525_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__nor2_4 _22166_ (.A(_05477_),
    .B(_05527_),
    .Y(_05528_));
 sky130_vsdinv _22167_ (.A(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hd__nand2_1 _22168_ (.A(_05527_),
    .B(_05477_),
    .Y(_05530_));
 sky130_fd_sc_hd__buf_6 _22169_ (.A(_14041_),
    .X(_05531_));
 sky130_fd_sc_hd__buf_6 _22170_ (.A(_05440_),
    .X(_05532_));
 sky130_fd_sc_hd__clkbuf_4 _22171_ (.A(_04716_),
    .X(_05533_));
 sky130_fd_sc_hd__nand3_2 _22172_ (.A(_05531_),
    .B(_05532_),
    .C(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hd__a22o_1 _22173_ (.A1(_14043_),
    .A2(_04719_),
    .B1(_05442_),
    .B2(_04874_),
    .X(_05535_));
 sky130_fd_sc_hd__o21a_1 _22174_ (.A1(_14449_),
    .A2(_05534_),
    .B1(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__and2_2 _22175_ (.A(_05355_),
    .B(_04928_),
    .X(_05537_));
 sky130_fd_sc_hd__nand2_2 _22176_ (.A(_14053_),
    .B(_04897_),
    .Y(_05538_));
 sky130_fd_sc_hd__and2_2 _22177_ (.A(_05357_),
    .B(_04988_),
    .X(_05539_));
 sky130_fd_sc_hd__xor2_4 _22178_ (.A(_05538_),
    .B(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__xor2_4 _22179_ (.A(_05537_),
    .B(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__xnor2_2 _22180_ (.A(_05536_),
    .B(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__a21oi_2 _22181_ (.A1(_05529_),
    .A2(_05530_),
    .B1(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__and3b_2 _22182_ (.A_N(_05528_),
    .B(_05542_),
    .C(_05530_),
    .X(_05544_));
 sky130_vsdinv _22183_ (.A(_05544_),
    .Y(_05545_));
 sky130_vsdinv _22184_ (.A(_05453_),
    .Y(_05546_));
 sky130_fd_sc_hd__nand3b_4 _22185_ (.A_N(_05543_),
    .B(_05545_),
    .C(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__o21bai_2 _22186_ (.A1(_05543_),
    .A2(_05544_),
    .B1_N(_05546_),
    .Y(_05548_));
 sky130_fd_sc_hd__nor2_2 _22187_ (.A(_05408_),
    .B(_05435_),
    .Y(_05549_));
 sky130_fd_sc_hd__a21oi_4 _22188_ (.A1(_05434_),
    .A2(_05410_),
    .B1(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__xor2_4 _22189_ (.A(_05550_),
    .B(_05438_),
    .X(_05551_));
 sky130_fd_sc_hd__a21oi_1 _22190_ (.A1(_05547_),
    .A2(_05548_),
    .B1(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__nand3_4 _22191_ (.A(_05547_),
    .B(_05548_),
    .C(_05551_),
    .Y(_05553_));
 sky130_vsdinv _22192_ (.A(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2_2 _22193_ (.A(_05461_),
    .B(_05456_),
    .Y(_05555_));
 sky130_fd_sc_hd__o21bai_2 _22194_ (.A1(_05552_),
    .A2(_05554_),
    .B1_N(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__a21o_1 _22195_ (.A1(_05547_),
    .A2(_05548_),
    .B1(_05551_),
    .X(_05557_));
 sky130_fd_sc_hd__nand3_4 _22196_ (.A(_05557_),
    .B(_05553_),
    .C(_05555_),
    .Y(_05558_));
 sky130_fd_sc_hd__and4_1 _22197_ (.A(_05351_),
    .B(_05348_),
    .C(_05350_),
    .D(_05458_),
    .X(_05559_));
 sky130_fd_sc_hd__a21oi_1 _22198_ (.A1(_05556_),
    .A2(_05558_),
    .B1(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand3_2 _22199_ (.A(_05556_),
    .B(_05559_),
    .C(_05558_),
    .Y(_05561_));
 sky130_vsdinv _22200_ (.A(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__a21o_1 _22201_ (.A1(_05468_),
    .A2(_05466_),
    .B1(_05465_),
    .X(_05563_));
 sky130_fd_sc_hd__o21bai_1 _22202_ (.A1(_05560_),
    .A2(_05562_),
    .B1_N(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__a21o_1 _22203_ (.A1(_05556_),
    .A2(_05558_),
    .B1(_05559_),
    .X(_05565_));
 sky130_fd_sc_hd__nand3_2 _22204_ (.A(_05565_),
    .B(_05561_),
    .C(_05563_),
    .Y(_05566_));
 sky130_fd_sc_hd__nand2_1 _22205_ (.A(_05564_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__a21oi_4 _22206_ (.A1(_05475_),
    .A2(_05474_),
    .B1(_05473_),
    .Y(_05568_));
 sky130_fd_sc_hd__xor2_1 _22207_ (.A(_05567_),
    .B(_05568_),
    .X(_02632_));
 sky130_fd_sc_hd__nand2_1 _22208_ (.A(_05553_),
    .B(_05547_),
    .Y(_05569_));
 sky130_fd_sc_hd__and2b_1 _22209_ (.A_N(_05480_),
    .B(_05492_),
    .X(_05570_));
 sky130_fd_sc_hd__o21bai_1 _22210_ (.A1(_05479_),
    .A2(_05493_),
    .B1_N(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__nor2_1 _22211_ (.A(_05489_),
    .B(_05490_),
    .Y(_05572_));
 sky130_fd_sc_hd__o21ba_1 _22212_ (.A1(_05482_),
    .A2(_05491_),
    .B1_N(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__or2b_4 _22213_ (.A(_05534_),
    .B_N(_04872_),
    .X(_05574_));
 sky130_fd_sc_hd__nand3b_4 _22214_ (.A_N(_05541_),
    .B(_05574_),
    .C(_05535_),
    .Y(_05575_));
 sky130_fd_sc_hd__clkbuf_4 _22215_ (.A(_14070_),
    .X(_05576_));
 sky130_fd_sc_hd__buf_2 _22216_ (.A(_05132_),
    .X(_05577_));
 sky130_fd_sc_hd__nand3b_1 _22217_ (.A_N(_05485_),
    .B(_05577_),
    .C(_05033_),
    .Y(_05578_));
 sky130_fd_sc_hd__o31a_4 _22218_ (.A1(_05576_),
    .A2(_14418_),
    .A3(_05488_),
    .B1(_05578_),
    .X(_05579_));
 sky130_fd_sc_hd__buf_6 _22219_ (.A(_14433_),
    .X(_05580_));
 sky130_fd_sc_hd__buf_4 _22220_ (.A(_14050_),
    .X(_05581_));
 sky130_fd_sc_hd__buf_6 _22221_ (.A(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__nand3b_1 _22222_ (.A_N(_05538_),
    .B(_05582_),
    .C(_04969_),
    .Y(_05583_));
 sky130_fd_sc_hd__o31a_2 _22223_ (.A1(_14059_),
    .A2(_05580_),
    .A3(_05540_),
    .B1(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__and2_2 _22224_ (.A(_05483_),
    .B(_05427_),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_4 _22225_ (.A(_14414_),
    .X(_05586_));
 sky130_fd_sc_hd__nand2_2 _22226_ (.A(_14066_),
    .B(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__buf_4 _22227_ (.A(_05129_),
    .X(_05588_));
 sky130_fd_sc_hd__and2_1 _22228_ (.A(_05588_),
    .B(_14420_),
    .X(_05589_));
 sky130_fd_sc_hd__xor2_4 _22229_ (.A(_05587_),
    .B(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__xor2_4 _22230_ (.A(_05585_),
    .B(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__xnor2_4 _22231_ (.A(_05584_),
    .B(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__xor2_4 _22232_ (.A(_05579_),
    .B(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__xor2_4 _22233_ (.A(_05575_),
    .B(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__xor2_2 _22234_ (.A(_05573_),
    .B(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__xnor2_1 _22235_ (.A(_05571_),
    .B(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__buf_6 _22236_ (.A(_05424_),
    .X(_05597_));
 sky130_fd_sc_hd__nor3_4 _22237_ (.A(_05302_),
    .B(_14401_),
    .C(_05507_),
    .Y(_05598_));
 sky130_fd_sc_hd__a41oi_4 _22238_ (.A1(_05299_),
    .A2(_04880_),
    .A3(_05597_),
    .A4(_05498_),
    .B1(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__nor2_1 _22239_ (.A(_05510_),
    .B(_05520_),
    .Y(_05600_));
 sky130_fd_sc_hd__o21bai_4 _22240_ (.A1(_05508_),
    .A2(_05521_),
    .B1_N(_05600_),
    .Y(_05601_));
 sky130_fd_sc_hd__and2_2 _22241_ (.A(_04933_),
    .B(_05498_),
    .X(_05602_));
 sky130_fd_sc_hd__nand2_2 _22242_ (.A(_04885_),
    .B(_05597_),
    .Y(_05603_));
 sky130_fd_sc_hd__buf_6 _22243_ (.A(_05513_),
    .X(_05604_));
 sky130_fd_sc_hd__nand2_2 _22244_ (.A(_04877_),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__xnor2_4 _22245_ (.A(_05603_),
    .B(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__xor2_4 _22246_ (.A(_05602_),
    .B(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__nand3b_1 _22247_ (.A_N(_05517_),
    .B(_05316_),
    .C(_05229_),
    .Y(_05608_));
 sky130_fd_sc_hd__o31a_2 _22248_ (.A1(_14098_),
    .A2(_14385_),
    .A3(_05519_),
    .B1(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__buf_4 _22249_ (.A(_14376_),
    .X(_05610_));
 sky130_fd_sc_hd__clkbuf_4 _22250_ (.A(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__and2_2 _22251_ (.A(_04714_),
    .B(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__clkbuf_4 _22252_ (.A(\pcpi_mul.rs1[10] ),
    .X(_05613_));
 sky130_fd_sc_hd__clkbuf_4 _22253_ (.A(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__nand2_2 _22254_ (.A(_05515_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__and2_2 _22255_ (.A(_05419_),
    .B(_05516_),
    .X(_05616_));
 sky130_fd_sc_hd__xor2_4 _22256_ (.A(_05615_),
    .B(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__xor2_4 _22257_ (.A(_05612_),
    .B(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__xnor2_4 _22258_ (.A(_05609_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__xor2_4 _22259_ (.A(_05607_),
    .B(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__xnor2_4 _22260_ (.A(_05601_),
    .B(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__xor2_4 _22261_ (.A(_05599_),
    .B(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__or2b_2 _22262_ (.A(_05596_),
    .B_N(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__or2b_2 _22263_ (.A(_05622_),
    .B_N(_05596_),
    .X(_05624_));
 sky130_fd_sc_hd__a21boi_1 _22264_ (.A1(_05495_),
    .A2(_05524_),
    .B1_N(_05496_),
    .Y(_05625_));
 sky130_fd_sc_hd__a21bo_1 _22265_ (.A1(_05623_),
    .A2(_05624_),
    .B1_N(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__nand3b_4 _22266_ (.A_N(_05625_),
    .B(_05623_),
    .C(_05624_),
    .Y(_05627_));
 sky130_fd_sc_hd__and2_1 _22267_ (.A(_05355_),
    .B(_05039_),
    .X(_05628_));
 sky130_fd_sc_hd__nand2_2 _22268_ (.A(_05447_),
    .B(_04956_),
    .Y(_05629_));
 sky130_fd_sc_hd__and2_2 _22269_ (.A(_14050_),
    .B(_04948_),
    .X(_05630_));
 sky130_fd_sc_hd__xor2_4 _22270_ (.A(_05629_),
    .B(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__xnor2_2 _22271_ (.A(_05628_),
    .B(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__nand2_4 _22272_ (.A(_05532_),
    .B(_04968_),
    .Y(_05633_));
 sky130_fd_sc_hd__clkbuf_2 _22273_ (.A(\pcpi_mul.rs2[14] ),
    .X(_05634_));
 sky130_fd_sc_hd__buf_4 _22274_ (.A(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__clkbuf_4 _22275_ (.A(\pcpi_mul.rs2[13] ),
    .X(_05636_));
 sky130_fd_sc_hd__buf_4 _22276_ (.A(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__nand3_4 _22277_ (.A(_05635_),
    .B(_05637_),
    .C(_04986_),
    .Y(_05638_));
 sky130_fd_sc_hd__a22o_1 _22278_ (.A1(_14036_),
    .A2(\pcpi_mul.rs1[0] ),
    .B1(_14041_),
    .B2(_04986_),
    .X(_05639_));
 sky130_fd_sc_hd__o21ai_4 _22279_ (.A1(_14451_),
    .A2(_05638_),
    .B1(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__xnor2_4 _22280_ (.A(_05633_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__xnor2_2 _22281_ (.A(_05574_),
    .B(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__xor2_2 _22282_ (.A(_05632_),
    .B(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__a21bo_1 _22283_ (.A1(_05626_),
    .A2(_05627_),
    .B1_N(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__nand3b_4 _22284_ (.A_N(_05643_),
    .B(_05626_),
    .C(_05627_),
    .Y(_05645_));
 sky130_fd_sc_hd__a21oi_1 _22285_ (.A1(_05644_),
    .A2(_05645_),
    .B1(_05544_),
    .Y(_05646_));
 sky130_fd_sc_hd__nor2_1 _22286_ (.A(_05500_),
    .B(_05523_),
    .Y(_05647_));
 sky130_fd_sc_hd__a21o_2 _22287_ (.A1(_05522_),
    .A2(_05502_),
    .B1(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__xor2_4 _22288_ (.A(_05648_),
    .B(_05528_),
    .X(_05649_));
 sky130_fd_sc_hd__nand3_4 _22289_ (.A(_05644_),
    .B(_05544_),
    .C(_05645_),
    .Y(_05650_));
 sky130_fd_sc_hd__nand3b_4 _22290_ (.A_N(_05646_),
    .B(_05649_),
    .C(_05650_),
    .Y(_05651_));
 sky130_vsdinv _22291_ (.A(_05650_),
    .Y(_05652_));
 sky130_fd_sc_hd__o21bai_1 _22292_ (.A1(_05646_),
    .A2(_05652_),
    .B1_N(_05649_),
    .Y(_05653_));
 sky130_fd_sc_hd__nand3_2 _22293_ (.A(_05569_),
    .B(_05651_),
    .C(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__a21o_1 _22294_ (.A1(_05653_),
    .A2(_05651_),
    .B1(_05569_),
    .X(_05655_));
 sky130_fd_sc_hd__o2bb2ai_1 _22295_ (.A1_N(_05654_),
    .A2_N(_05655_),
    .B1(_05438_),
    .B2(_05550_),
    .Y(_05656_));
 sky130_fd_sc_hd__a211oi_4 _22296_ (.A1(_05348_),
    .A2(_05387_),
    .B1(_05550_),
    .C1(_05437_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand3_2 _22297_ (.A(_05655_),
    .B(_05657_),
    .C(_05654_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2_1 _22298_ (.A(_05561_),
    .B(_05558_),
    .Y(_05659_));
 sky130_fd_sc_hd__a21oi_2 _22299_ (.A1(_05656_),
    .A2(_05658_),
    .B1(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__and3_2 _22300_ (.A(_05656_),
    .B(_05659_),
    .C(_05658_),
    .X(_05661_));
 sky130_fd_sc_hd__nor2_4 _22301_ (.A(_05660_),
    .B(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__o21ai_2 _22302_ (.A1(_05567_),
    .A2(_05568_),
    .B1(_05566_),
    .Y(_05663_));
 sky130_fd_sc_hd__xor2_1 _22303_ (.A(_05662_),
    .B(_05663_),
    .X(_02633_));
 sky130_fd_sc_hd__nand3b_1 _22304_ (.A_N(_05541_),
    .B(_05593_),
    .C(_05536_),
    .Y(_05664_));
 sky130_fd_sc_hd__o21a_1 _22305_ (.A1(_05573_),
    .A2(_05594_),
    .B1(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__nor2_1 _22306_ (.A(_05584_),
    .B(_05591_),
    .Y(_05666_));
 sky130_fd_sc_hd__o21ba_2 _22307_ (.A1(_05579_),
    .A2(_05592_),
    .B1_N(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__or2b_1 _22308_ (.A(_05642_),
    .B_N(_05632_),
    .X(_05668_));
 sky130_fd_sc_hd__o21ai_4 _22309_ (.A1(_05574_),
    .A2(_05641_),
    .B1(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__nand3b_2 _22310_ (.A_N(_05587_),
    .B(_05337_),
    .C(_05092_),
    .Y(_05670_));
 sky130_fd_sc_hd__o31a_4 _22311_ (.A1(_14071_),
    .A2(_14412_),
    .A3(_05590_),
    .B1(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__nand3b_1 _22312_ (.A_N(_05629_),
    .B(_05582_),
    .C(_04974_),
    .Y(_05672_));
 sky130_fd_sc_hd__o31a_2 _22313_ (.A1(_14059_),
    .A2(_05247_),
    .A3(_05631_),
    .B1(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__and2_2 _22314_ (.A(_04997_),
    .B(_05308_),
    .X(_05674_));
 sky130_fd_sc_hd__nand2_2 _22315_ (.A(_05163_),
    .B(_05227_),
    .Y(_05675_));
 sky130_fd_sc_hd__and2_1 _22316_ (.A(_05486_),
    .B(_05586_),
    .X(_05676_));
 sky130_fd_sc_hd__xor2_4 _22317_ (.A(_05675_),
    .B(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__xor2_4 _22318_ (.A(_05674_),
    .B(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__xnor2_4 _22319_ (.A(_05673_),
    .B(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__xor2_4 _22320_ (.A(_05671_),
    .B(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__xnor2_4 _22321_ (.A(_05669_),
    .B(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__xor2_4 _22322_ (.A(_05667_),
    .B(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__xor2_2 _22323_ (.A(_05665_),
    .B(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__nor3_4 _22324_ (.A(_05302_),
    .B(_14395_),
    .C(_05606_),
    .Y(_05684_));
 sky130_fd_sc_hd__a41oi_4 _22325_ (.A1(_05299_),
    .A2(_04880_),
    .A3(_05604_),
    .A4(_05597_),
    .B1(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__nor2_1 _22326_ (.A(_05609_),
    .B(_05618_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21bai_4 _22327_ (.A1(_05607_),
    .A2(_05619_),
    .B1_N(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__and2_2 _22328_ (.A(_04933_),
    .B(_05597_),
    .X(_05688_));
 sky130_fd_sc_hd__nand2_2 _22329_ (.A(_04885_),
    .B(_05604_),
    .Y(_05689_));
 sky130_fd_sc_hd__buf_2 _22330_ (.A(_14376_),
    .X(_05690_));
 sky130_fd_sc_hd__clkbuf_4 _22331_ (.A(_05690_),
    .X(_05691_));
 sky130_fd_sc_hd__buf_6 _22332_ (.A(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_2 _22333_ (.A(_04877_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__xnor2_4 _22334_ (.A(_05689_),
    .B(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__xor2_4 _22335_ (.A(_05688_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__nand3b_1 _22336_ (.A_N(_05615_),
    .B(_05316_),
    .C(_05301_),
    .Y(_05696_));
 sky130_fd_sc_hd__o31a_2 _22337_ (.A1(_14098_),
    .A2(_14379_),
    .A3(_05617_),
    .B1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__buf_2 _22338_ (.A(\pcpi_mul.rs1[15] ),
    .X(_05698_));
 sky130_fd_sc_hd__buf_6 _22339_ (.A(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__clkbuf_4 _22340_ (.A(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__and2_2 _22341_ (.A(_04714_),
    .B(_05700_),
    .X(_05701_));
 sky130_fd_sc_hd__nand2_2 _22342_ (.A(_05515_),
    .B(_05497_),
    .Y(_05702_));
 sky130_fd_sc_hd__and2_1 _22343_ (.A(_05419_),
    .B(_05241_),
    .X(_05703_));
 sky130_fd_sc_hd__xor2_4 _22344_ (.A(_05702_),
    .B(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__xor2_4 _22345_ (.A(_05701_),
    .B(_05704_),
    .X(_05705_));
 sky130_fd_sc_hd__xnor2_4 _22346_ (.A(_05697_),
    .B(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__xor2_4 _22347_ (.A(_05695_),
    .B(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__xnor2_4 _22348_ (.A(_05687_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__xor2_4 _22349_ (.A(_05685_),
    .B(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__nand2b_4 _22350_ (.A_N(_05683_),
    .B(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__or2b_2 _22351_ (.A(_05709_),
    .B_N(_05683_),
    .X(_05711_));
 sky130_fd_sc_hd__nand2_1 _22352_ (.A(_05595_),
    .B(_05571_),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_2 _22353_ (.A(_05623_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__a21o_1 _22354_ (.A1(_05710_),
    .A2(_05711_),
    .B1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__nand3_4 _22355_ (.A(_05713_),
    .B(_05710_),
    .C(_05711_),
    .Y(_05715_));
 sky130_fd_sc_hd__clkbuf_4 _22356_ (.A(\pcpi_mul.rs2[15] ),
    .X(_05716_));
 sky130_fd_sc_hd__clkbuf_4 _22357_ (.A(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__clkbuf_4 _22358_ (.A(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__and2_2 _22359_ (.A(net438),
    .B(_04720_),
    .X(_05719_));
 sky130_fd_sc_hd__buf_4 _22360_ (.A(_05354_),
    .X(_05720_));
 sky130_fd_sc_hd__and2_2 _22361_ (.A(_05720_),
    .B(_05092_),
    .X(_05721_));
 sky130_fd_sc_hd__nand2_2 _22362_ (.A(_05447_),
    .B(_04960_),
    .Y(_05722_));
 sky130_fd_sc_hd__and2_1 _22363_ (.A(_05357_),
    .B(_14432_),
    .X(_05723_));
 sky130_fd_sc_hd__xor2_4 _22364_ (.A(_05722_),
    .B(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__xnor2_4 _22365_ (.A(_05721_),
    .B(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__o22a_4 _22366_ (.A1(_14452_),
    .A2(_05638_),
    .B1(_05633_),
    .B2(_05640_),
    .X(_05726_));
 sky130_fd_sc_hd__buf_4 _22367_ (.A(\pcpi_mul.rs2[12] ),
    .X(_05727_));
 sky130_fd_sc_hd__buf_4 _22368_ (.A(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__and2_2 _22369_ (.A(_05728_),
    .B(_05051_),
    .X(_05729_));
 sky130_fd_sc_hd__buf_4 _22370_ (.A(\pcpi_mul.rs2[14] ),
    .X(_05730_));
 sky130_fd_sc_hd__nand2_2 _22371_ (.A(_05730_),
    .B(_14447_),
    .Y(_05731_));
 sky130_fd_sc_hd__buf_4 _22372_ (.A(_05636_),
    .X(_05732_));
 sky130_fd_sc_hd__nand2_2 _22373_ (.A(_05732_),
    .B(_04988_),
    .Y(_05733_));
 sky130_fd_sc_hd__xnor2_4 _22374_ (.A(_05731_),
    .B(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__xor2_4 _22375_ (.A(_05729_),
    .B(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__xnor2_4 _22376_ (.A(_05726_),
    .B(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__xnor2_4 _22377_ (.A(_05725_),
    .B(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__xor2_4 _22378_ (.A(_05719_),
    .B(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__a21o_1 _22379_ (.A1(_05714_),
    .A2(_05715_),
    .B1(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__nand3_4 _22380_ (.A(_05714_),
    .B(_05738_),
    .C(_05715_),
    .Y(_05740_));
 sky130_vsdinv _22381_ (.A(_05645_),
    .Y(_05741_));
 sky130_fd_sc_hd__a21oi_4 _22382_ (.A1(_05739_),
    .A2(_05740_),
    .B1(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__nand3_4 _22383_ (.A(_05739_),
    .B(_05741_),
    .C(_05740_),
    .Y(_05743_));
 sky130_vsdinv _22384_ (.A(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__nor2_2 _22385_ (.A(_05599_),
    .B(_05621_),
    .Y(_05745_));
 sky130_fd_sc_hd__a21oi_4 _22386_ (.A1(_05620_),
    .A2(_05601_),
    .B1(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__xor2_4 _22387_ (.A(_05746_),
    .B(_05627_),
    .X(_05747_));
 sky130_fd_sc_hd__o21bai_2 _22388_ (.A1(_05742_),
    .A2(_05744_),
    .B1_N(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand3b_4 _22389_ (.A_N(_05742_),
    .B(_05747_),
    .C(_05743_),
    .Y(_05749_));
 sky130_fd_sc_hd__nand2_2 _22390_ (.A(_05651_),
    .B(_05650_),
    .Y(_05750_));
 sky130_fd_sc_hd__a21o_1 _22391_ (.A1(_05748_),
    .A2(_05749_),
    .B1(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__nand3_4 _22392_ (.A(_05750_),
    .B(_05749_),
    .C(_05748_),
    .Y(_05752_));
 sky130_fd_sc_hd__nor3b_4 _22393_ (.A(_05477_),
    .B(_05527_),
    .C_N(_05648_),
    .Y(_05753_));
 sky130_fd_sc_hd__a21o_1 _22394_ (.A1(_05751_),
    .A2(_05752_),
    .B1(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__nand3_4 _22395_ (.A(_05751_),
    .B(_05753_),
    .C(_05752_),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _22396_ (.A(_05658_),
    .B(_05654_),
    .Y(_05756_));
 sky130_fd_sc_hd__a21oi_1 _22397_ (.A1(_05754_),
    .A2(_05755_),
    .B1(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__and3_1 _22398_ (.A(_05754_),
    .B(_05756_),
    .C(_05755_),
    .X(_05758_));
 sky130_fd_sc_hd__nor2_1 _22399_ (.A(_05757_),
    .B(_05758_),
    .Y(_05759_));
 sky130_vsdinv _22400_ (.A(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__a21oi_4 _22401_ (.A1(_05663_),
    .A2(_05662_),
    .B1(_05661_),
    .Y(_05761_));
 sky130_fd_sc_hd__xor2_1 _22402_ (.A(_05760_),
    .B(_05761_),
    .X(_02634_));
 sky130_fd_sc_hd__nor3_4 _22403_ (.A(_05302_),
    .B(_14390_),
    .C(_05694_),
    .Y(_05762_));
 sky130_fd_sc_hd__a41oi_4 _22404_ (.A1(_05299_),
    .A2(_04880_),
    .A3(_05692_),
    .A4(_05604_),
    .B1(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__nor2_1 _22405_ (.A(_05697_),
    .B(_05705_),
    .Y(_05764_));
 sky130_fd_sc_hd__o21bai_4 _22406_ (.A1(_05695_),
    .A2(_05706_),
    .B1_N(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__and2_2 _22407_ (.A(_04933_),
    .B(_05604_),
    .X(_05766_));
 sky130_fd_sc_hd__nand2_2 _22408_ (.A(_04905_),
    .B(_05692_),
    .Y(_05767_));
 sky130_fd_sc_hd__clkbuf_4 _22409_ (.A(_14370_),
    .X(_05768_));
 sky130_fd_sc_hd__clkbuf_4 _22410_ (.A(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__buf_4 _22411_ (.A(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__nand2_2 _22412_ (.A(_04877_),
    .B(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__xnor2_4 _22413_ (.A(_05767_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__xor2_4 _22414_ (.A(_05766_),
    .B(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__nand3b_1 _22415_ (.A_N(_05702_),
    .B(_05316_),
    .C(_05406_),
    .Y(_05774_));
 sky130_fd_sc_hd__o31a_2 _22416_ (.A1(_14098_),
    .A2(_14373_),
    .A3(_05704_),
    .B1(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__clkbuf_4 _22417_ (.A(\pcpi_mul.rs1[16] ),
    .X(_05776_));
 sky130_fd_sc_hd__clkbuf_4 _22418_ (.A(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__clkbuf_4 _22419_ (.A(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__and2_2 _22420_ (.A(_04714_),
    .B(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__nand2_2 _22421_ (.A(_05324_),
    .B(_05423_),
    .Y(_05780_));
 sky130_fd_sc_hd__and2_1 _22422_ (.A(_05326_),
    .B(_05321_),
    .X(_05781_));
 sky130_fd_sc_hd__xor2_4 _22423_ (.A(_05780_),
    .B(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__xor2_4 _22424_ (.A(_05779_),
    .B(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__xnor2_4 _22425_ (.A(_05775_),
    .B(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__xor2_4 _22426_ (.A(_05773_),
    .B(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__xnor2_4 _22427_ (.A(_05765_),
    .B(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__xor2_4 _22428_ (.A(_05763_),
    .B(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__and2_1 _22429_ (.A(_05680_),
    .B(_05669_),
    .X(_05788_));
 sky130_fd_sc_hd__o21ba_1 _22430_ (.A1(_05667_),
    .A2(_05681_),
    .B1_N(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__nor2_1 _22431_ (.A(_05673_),
    .B(_05678_),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ba_2 _22432_ (.A1(_05671_),
    .A2(_05679_),
    .B1_N(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__or2b_1 _22433_ (.A(_05736_),
    .B_N(_05725_),
    .X(_05792_));
 sky130_fd_sc_hd__o21ai_4 _22434_ (.A1(_05735_),
    .A2(_05726_),
    .B1(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__nand3b_1 _22435_ (.A_N(_05675_),
    .B(_05337_),
    .C(_05191_),
    .Y(_05794_));
 sky130_fd_sc_hd__o31a_4 _22436_ (.A1(_05576_),
    .A2(_14406_),
    .A3(_05677_),
    .B1(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__nand3b_1 _22437_ (.A_N(_05722_),
    .B(_05582_),
    .C(_04928_),
    .Y(_05796_));
 sky130_fd_sc_hd__o31a_2 _22438_ (.A1(_14059_),
    .A2(_05057_),
    .A3(_05724_),
    .B1(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__and2_2 _22439_ (.A(_05483_),
    .B(_05241_),
    .X(_05798_));
 sky130_fd_sc_hd__nand2_2 _22440_ (.A(_14066_),
    .B(_05236_),
    .Y(_05799_));
 sky130_fd_sc_hd__and2_1 _22441_ (.A(_05588_),
    .B(_05426_),
    .X(_05800_));
 sky130_fd_sc_hd__xor2_4 _22442_ (.A(_05799_),
    .B(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__xor2_4 _22443_ (.A(_05798_),
    .B(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__xnor2_4 _22444_ (.A(_05797_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__xor2_4 _22445_ (.A(_05795_),
    .B(_05803_),
    .X(_05804_));
 sky130_fd_sc_hd__xnor2_4 _22446_ (.A(_05793_),
    .B(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__xor2_4 _22447_ (.A(_05791_),
    .B(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__xnor2_2 _22448_ (.A(_05789_),
    .B(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__xor2_4 _22449_ (.A(_05787_),
    .B(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__or2b_2 _22450_ (.A(_05665_),
    .B_N(_05682_),
    .X(_05809_));
 sky130_fd_sc_hd__nand2_2 _22451_ (.A(_05710_),
    .B(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand2_8 _22452_ (.A(_05808_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__nand3b_4 _22453_ (.A_N(_05808_),
    .B(_05809_),
    .C(_05710_),
    .Y(_05812_));
 sky130_fd_sc_hd__nand2_2 _22454_ (.A(_05737_),
    .B(_05719_),
    .Y(_05813_));
 sky130_fd_sc_hd__clkbuf_8 _22455_ (.A(_14027_),
    .X(_05814_));
 sky130_fd_sc_hd__clkbuf_8 _22456_ (.A(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__nand2_4 _22457_ (.A(_05815_),
    .B(_04718_),
    .Y(_05816_));
 sky130_fd_sc_hd__nand2_4 _22458_ (.A(net438),
    .B(_04873_),
    .Y(_05817_));
 sky130_fd_sc_hd__xor2_4 _22459_ (.A(_05816_),
    .B(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__buf_4 _22460_ (.A(_05048_),
    .X(_05819_));
 sky130_fd_sc_hd__and2_2 _22461_ (.A(_05720_),
    .B(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__nand2_2 _22462_ (.A(_05271_),
    .B(_05090_),
    .Y(_05821_));
 sky130_fd_sc_hd__and2_1 _22463_ (.A(\pcpi_mul.rs2[11] ),
    .B(_04959_),
    .X(_05822_));
 sky130_fd_sc_hd__xor2_4 _22464_ (.A(_05821_),
    .B(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__xor2_4 _22465_ (.A(_05820_),
    .B(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__and2_2 _22466_ (.A(_05728_),
    .B(_04927_),
    .X(_05825_));
 sky130_fd_sc_hd__nand2_2 _22467_ (.A(_14041_),
    .B(_04948_),
    .Y(_05826_));
 sky130_fd_sc_hd__and2_1 _22468_ (.A(_05730_),
    .B(_14441_),
    .X(_05827_));
 sky130_fd_sc_hd__xor2_4 _22469_ (.A(_05826_),
    .B(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__xor2_4 _22470_ (.A(_05825_),
    .B(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__o32a_4 _22471_ (.A1(_14047_),
    .A2(_14438_),
    .A3(_05734_),
    .B1(_14443_),
    .B2(_05638_),
    .X(_05830_));
 sky130_fd_sc_hd__xnor2_4 _22472_ (.A(_05829_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__xor2_4 _22473_ (.A(_05824_),
    .B(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__xnor2_4 _22474_ (.A(_05818_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__nor2_4 _22475_ (.A(_05813_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__and2_1 _22476_ (.A(_05833_),
    .B(_05813_),
    .X(_05835_));
 sky130_fd_sc_hd__o2bb2ai_4 _22477_ (.A1_N(_05811_),
    .A2_N(_05812_),
    .B1(_05834_),
    .B2(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__xor2_2 _22478_ (.A(_05813_),
    .B(_05833_),
    .X(_05837_));
 sky130_fd_sc_hd__nand3_4 _22479_ (.A(_05812_),
    .B(_05837_),
    .C(_05811_),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2_4 _22480_ (.A(_05836_),
    .B(_05838_),
    .Y(_05839_));
 sky130_fd_sc_hd__nand2_2 _22481_ (.A(_05839_),
    .B(_05740_),
    .Y(_05840_));
 sky130_vsdinv _22482_ (.A(_05740_),
    .Y(_05841_));
 sky130_fd_sc_hd__nand3_2 _22483_ (.A(_05841_),
    .B(_05836_),
    .C(_05838_),
    .Y(_05842_));
 sky130_fd_sc_hd__nor2_2 _22484_ (.A(_05685_),
    .B(_05708_),
    .Y(_05843_));
 sky130_fd_sc_hd__a21oi_4 _22485_ (.A1(_05707_),
    .A2(_05687_),
    .B1(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__xor2_4 _22486_ (.A(_05844_),
    .B(_05715_),
    .X(_05845_));
 sky130_fd_sc_hd__a21oi_1 _22487_ (.A1(_05840_),
    .A2(_05842_),
    .B1(_05845_),
    .Y(_05846_));
 sky130_vsdinv _22488_ (.A(_05845_),
    .Y(_05847_));
 sky130_fd_sc_hd__a21oi_4 _22489_ (.A1(_05836_),
    .A2(_05838_),
    .B1(_05841_),
    .Y(_05848_));
 sky130_fd_sc_hd__nor2_8 _22490_ (.A(_05740_),
    .B(_05839_),
    .Y(_05849_));
 sky130_fd_sc_hd__nor3_4 _22491_ (.A(_05847_),
    .B(_05848_),
    .C(_05849_),
    .Y(_05850_));
 sky130_vsdinv _22492_ (.A(_05747_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21ai_2 _22493_ (.A1(_05851_),
    .A2(_05742_),
    .B1(_05743_),
    .Y(_05852_));
 sky130_fd_sc_hd__o21bai_2 _22494_ (.A1(_05846_),
    .A2(_05850_),
    .B1_N(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__o21bai_2 _22495_ (.A1(_05848_),
    .A2(_05849_),
    .B1_N(_05845_),
    .Y(_05854_));
 sky130_fd_sc_hd__nand3_2 _22496_ (.A(_05840_),
    .B(_05845_),
    .C(_05842_),
    .Y(_05855_));
 sky130_fd_sc_hd__nand3_4 _22497_ (.A(_05854_),
    .B(_05855_),
    .C(_05852_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_1 _22498_ (.A(_05853_),
    .B(_05856_),
    .Y(_05857_));
 sky130_fd_sc_hd__nor2_4 _22499_ (.A(_05746_),
    .B(_05627_),
    .Y(_05858_));
 sky130_vsdinv _22500_ (.A(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__nand2_2 _22501_ (.A(_05857_),
    .B(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__nand3_4 _22502_ (.A(_05853_),
    .B(_05858_),
    .C(_05856_),
    .Y(_05861_));
 sky130_fd_sc_hd__nand2_1 _22503_ (.A(_05755_),
    .B(_05752_),
    .Y(_05862_));
 sky130_fd_sc_hd__a21oi_2 _22504_ (.A1(_05860_),
    .A2(_05861_),
    .B1(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__nand2_1 _22505_ (.A(_05860_),
    .B(_05861_),
    .Y(_05864_));
 sky130_fd_sc_hd__a21oi_4 _22506_ (.A1(_05752_),
    .A2(_05755_),
    .B1(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__nor2_4 _22507_ (.A(_05863_),
    .B(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__o21bai_4 _22508_ (.A1(_05760_),
    .A2(_05761_),
    .B1_N(_05758_),
    .Y(_05867_));
 sky130_fd_sc_hd__buf_4 _22509_ (.A(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__xor2_1 _22510_ (.A(_05866_),
    .B(_05868_),
    .X(_02635_));
 sky130_fd_sc_hd__a21oi_4 _22511_ (.A1(_05840_),
    .A2(_05845_),
    .B1(_05849_),
    .Y(_05869_));
 sky130_fd_sc_hd__nor2_1 _22512_ (.A(_05797_),
    .B(_05802_),
    .Y(_05870_));
 sky130_fd_sc_hd__nor2_1 _22513_ (.A(_05795_),
    .B(_05803_),
    .Y(_05871_));
 sky130_fd_sc_hd__nor2_1 _22514_ (.A(_05829_),
    .B(_05830_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21bai_2 _22515_ (.A1(_05824_),
    .A2(_05831_),
    .B1_N(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__buf_6 _22516_ (.A(_14399_),
    .X(_05874_));
 sky130_fd_sc_hd__buf_4 _22517_ (.A(_05106_),
    .X(_05875_));
 sky130_fd_sc_hd__nand3b_1 _22518_ (.A_N(_05799_),
    .B(_05127_),
    .C(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__o31a_4 _22519_ (.A1(_14070_),
    .A2(_05874_),
    .A3(_05801_),
    .B1(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__buf_4 _22520_ (.A(_14058_),
    .X(_05878_));
 sky130_fd_sc_hd__buf_6 _22521_ (.A(_05445_),
    .X(_05879_));
 sky130_fd_sc_hd__nand3b_2 _22522_ (.A_N(_05821_),
    .B(_05879_),
    .C(_05032_),
    .Y(_05880_));
 sky130_fd_sc_hd__o31a_4 _22523_ (.A1(_05878_),
    .A2(_14417_),
    .A3(_05823_),
    .B1(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__clkbuf_4 _22524_ (.A(\pcpi_mul.rs1[11] ),
    .X(_05882_));
 sky130_fd_sc_hd__and2_2 _22525_ (.A(_04996_),
    .B(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__clkbuf_4 _22526_ (.A(_14065_),
    .X(_05884_));
 sky130_fd_sc_hd__nand2_2 _22527_ (.A(_05884_),
    .B(_14398_),
    .Y(_05885_));
 sky130_fd_sc_hd__and2_1 _22528_ (.A(_14061_),
    .B(\pcpi_mul.rs1[9] ),
    .X(_05886_));
 sky130_fd_sc_hd__xor2_4 _22529_ (.A(_05885_),
    .B(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__xor2_4 _22530_ (.A(_05883_),
    .B(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__xnor2_4 _22531_ (.A(_05881_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__xor2_4 _22532_ (.A(_05877_),
    .B(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__xnor2_1 _22533_ (.A(_05873_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__o21bai_2 _22534_ (.A1(_05870_),
    .A2(_05871_),
    .B1_N(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__o21ba_1 _22535_ (.A1(_05795_),
    .A2(_05803_),
    .B1_N(_05870_),
    .X(_05893_));
 sky130_fd_sc_hd__nand2_2 _22536_ (.A(_05891_),
    .B(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__and2_1 _22537_ (.A(_05804_),
    .B(_05793_),
    .X(_05895_));
 sky130_fd_sc_hd__o21bai_2 _22538_ (.A1(_05791_),
    .A2(_05805_),
    .B1_N(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__a21oi_4 _22539_ (.A1(_05892_),
    .A2(_05894_),
    .B1(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__and3_2 _22540_ (.A(_05892_),
    .B(_05896_),
    .C(_05894_),
    .X(_05898_));
 sky130_fd_sc_hd__buf_6 _22541_ (.A(_04878_),
    .X(_05899_));
 sky130_fd_sc_hd__nand3b_2 _22542_ (.A_N(_05767_),
    .B(_05899_),
    .C(_05770_),
    .Y(_05900_));
 sky130_fd_sc_hd__o31ai_4 _22543_ (.A1(_14088_),
    .A2(_14385_),
    .A3(_05772_),
    .B1(_05900_),
    .Y(_05901_));
 sky130_fd_sc_hd__nor2_1 _22544_ (.A(_05775_),
    .B(_05783_),
    .Y(_05902_));
 sky130_fd_sc_hd__o21bai_4 _22545_ (.A1(_05773_),
    .A2(_05784_),
    .B1_N(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__and2_2 _22546_ (.A(_14083_),
    .B(_05692_),
    .X(_05904_));
 sky130_fd_sc_hd__clkbuf_4 _22547_ (.A(_05768_),
    .X(_05905_));
 sky130_fd_sc_hd__nand2_2 _22548_ (.A(_04936_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__nand2_2 _22549_ (.A(_04938_),
    .B(_05778_),
    .Y(_05907_));
 sky130_fd_sc_hd__xnor2_4 _22550_ (.A(_05906_),
    .B(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__xor2_4 _22551_ (.A(_05904_),
    .B(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__nand3b_1 _22552_ (.A_N(_05780_),
    .B(_05420_),
    .C(_05498_),
    .Y(_05910_));
 sky130_fd_sc_hd__o31a_2 _22553_ (.A1(_05315_),
    .A2(_14367_),
    .A3(_05782_),
    .B1(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__buf_6 _22554_ (.A(_14357_),
    .X(_05912_));
 sky130_fd_sc_hd__clkbuf_4 _22555_ (.A(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__and2_2 _22556_ (.A(_04955_),
    .B(_05913_),
    .X(_05914_));
 sky130_fd_sc_hd__buf_2 _22557_ (.A(_14381_),
    .X(_05915_));
 sky130_fd_sc_hd__nand2_2 _22558_ (.A(_04924_),
    .B(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__clkbuf_4 _22559_ (.A(\pcpi_mul.rs1[12] ),
    .X(_05917_));
 sky130_fd_sc_hd__and2_1 _22560_ (.A(_14073_),
    .B(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__xor2_4 _22561_ (.A(_05916_),
    .B(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__xor2_4 _22562_ (.A(_05914_),
    .B(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__xnor2_4 _22563_ (.A(_05911_),
    .B(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__xor2_4 _22564_ (.A(_05909_),
    .B(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__xnor2_4 _22565_ (.A(_05903_),
    .B(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__xnor2_4 _22566_ (.A(_05901_),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__nor3b_4 _22567_ (.A(_05897_),
    .B(_05898_),
    .C_N(_05924_),
    .Y(_05925_));
 sky130_fd_sc_hd__o21ba_1 _22568_ (.A1(_05897_),
    .A2(_05898_),
    .B1_N(_05924_),
    .X(_05926_));
 sky130_fd_sc_hd__nor3b_4 _22569_ (.A(_05925_),
    .B(_05926_),
    .C_N(_05834_),
    .Y(_05927_));
 sky130_fd_sc_hd__o21bai_2 _22570_ (.A1(_05925_),
    .A2(_05926_),
    .B1_N(_05834_),
    .Y(_05928_));
 sky130_vsdinv _22571_ (.A(_05928_),
    .Y(_05929_));
 sky130_fd_sc_hd__or2b_1 _22572_ (.A(_05806_),
    .B_N(_05789_),
    .X(_05930_));
 sky130_fd_sc_hd__and2b_1 _22573_ (.A_N(_05789_),
    .B(_05806_),
    .X(_05931_));
 sky130_fd_sc_hd__a21oi_1 _22574_ (.A1(_05930_),
    .A2(_05787_),
    .B1(_05931_),
    .Y(_05932_));
 sky130_vsdinv _22575_ (.A(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__o21bai_2 _22576_ (.A1(_05927_),
    .A2(_05929_),
    .B1_N(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__nand3b_4 _22577_ (.A_N(_05927_),
    .B(_05933_),
    .C(_05928_),
    .Y(_05935_));
 sky130_fd_sc_hd__nand2_2 _22578_ (.A(_05934_),
    .B(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__nand2_4 _22579_ (.A(_05832_),
    .B(_05818_),
    .Y(_05937_));
 sky130_fd_sc_hd__nor2_4 _22580_ (.A(_05816_),
    .B(_05817_),
    .Y(_05938_));
 sky130_fd_sc_hd__buf_6 _22581_ (.A(_05716_),
    .X(_05939_));
 sky130_fd_sc_hd__nand2_2 _22582_ (.A(_05939_),
    .B(_04937_),
    .Y(_05940_));
 sky130_fd_sc_hd__buf_6 _22583_ (.A(_14023_),
    .X(_05941_));
 sky130_fd_sc_hd__nand3_4 _22584_ (.A(_05941_),
    .B(_05814_),
    .C(_04907_),
    .Y(_05942_));
 sky130_fd_sc_hd__buf_4 _22585_ (.A(_14023_),
    .X(_05943_));
 sky130_fd_sc_hd__buf_4 _22586_ (.A(_14027_),
    .X(_05944_));
 sky130_fd_sc_hd__a22o_1 _22587_ (.A1(_05943_),
    .A2(_05533_),
    .B1(_05944_),
    .B2(_04907_),
    .X(_05945_));
 sky130_fd_sc_hd__o21ai_4 _22588_ (.A1(_14453_),
    .A2(_05942_),
    .B1(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__xnor2_4 _22589_ (.A(_05940_),
    .B(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__xnor2_4 _22590_ (.A(_05938_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__and2_2 _22591_ (.A(_05720_),
    .B(_05875_),
    .X(_05949_));
 sky130_fd_sc_hd__nand2_2 _22592_ (.A(_05271_),
    .B(_05046_),
    .Y(_05950_));
 sky130_fd_sc_hd__and2_1 _22593_ (.A(\pcpi_mul.rs2[11] ),
    .B(_05089_),
    .X(_05951_));
 sky130_fd_sc_hd__xor2_4 _22594_ (.A(_05950_),
    .B(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__xor2_4 _22595_ (.A(_05949_),
    .B(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__buf_4 _22596_ (.A(\pcpi_mul.rs2[14] ),
    .X(_05954_));
 sky130_fd_sc_hd__clkbuf_4 _22597_ (.A(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__buf_6 _22598_ (.A(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__nand3b_1 _22599_ (.A_N(_05826_),
    .B(_05956_),
    .C(_04969_),
    .Y(_05957_));
 sky130_fd_sc_hd__o31a_2 _22600_ (.A1(_14047_),
    .A2(_05580_),
    .A3(_05828_),
    .B1(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__clkbuf_4 _22601_ (.A(_14426_),
    .X(_05959_));
 sky130_fd_sc_hd__and2_2 _22602_ (.A(_05728_),
    .B(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__nand2_2 _22603_ (.A(_05637_),
    .B(_14432_),
    .Y(_05961_));
 sky130_fd_sc_hd__and2_1 _22604_ (.A(_05730_),
    .B(_04948_),
    .X(_05962_));
 sky130_fd_sc_hd__xor2_4 _22605_ (.A(_05961_),
    .B(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__xor2_4 _22606_ (.A(_05960_),
    .B(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__xnor2_4 _22607_ (.A(_05958_),
    .B(_05964_),
    .Y(_05965_));
 sky130_fd_sc_hd__xor2_4 _22608_ (.A(_05953_),
    .B(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__xnor2_4 _22609_ (.A(_05948_),
    .B(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__xor2_4 _22610_ (.A(_05937_),
    .B(_05967_),
    .X(_05968_));
 sky130_vsdinv _22611_ (.A(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand2_2 _22612_ (.A(_05936_),
    .B(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__nand3_4 _22613_ (.A(_05934_),
    .B(_05968_),
    .C(_05935_),
    .Y(_05971_));
 sky130_vsdinv _22614_ (.A(_05838_),
    .Y(_05972_));
 sky130_fd_sc_hd__a21o_1 _22615_ (.A1(_05970_),
    .A2(_05971_),
    .B1(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__nand3_4 _22616_ (.A(_05972_),
    .B(_05970_),
    .C(_05971_),
    .Y(_05974_));
 sky130_fd_sc_hd__nor2_2 _22617_ (.A(_05763_),
    .B(_05786_),
    .Y(_05975_));
 sky130_fd_sc_hd__a21oi_4 _22618_ (.A1(_05785_),
    .A2(_05765_),
    .B1(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__xor2_4 _22619_ (.A(_05976_),
    .B(_05811_),
    .X(_05977_));
 sky130_fd_sc_hd__a21o_1 _22620_ (.A1(_05973_),
    .A2(_05974_),
    .B1(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__nand3_4 _22621_ (.A(_05973_),
    .B(_05977_),
    .C(_05974_),
    .Y(_05979_));
 sky130_fd_sc_hd__nand3b_4 _22622_ (.A_N(_05869_),
    .B(_05978_),
    .C(_05979_),
    .Y(_05980_));
 sky130_fd_sc_hd__a21oi_2 _22623_ (.A1(_05973_),
    .A2(_05974_),
    .B1(_05977_),
    .Y(_05981_));
 sky130_vsdinv _22624_ (.A(_05979_),
    .Y(_05982_));
 sky130_fd_sc_hd__o21ai_4 _22625_ (.A1(_05981_),
    .A2(_05982_),
    .B1(_05869_),
    .Y(_05983_));
 sky130_fd_sc_hd__o2bb2ai_4 _22626_ (.A1_N(_05980_),
    .A2_N(_05983_),
    .B1(_05715_),
    .B2(_05844_),
    .Y(_05984_));
 sky130_fd_sc_hd__nor2_2 _22627_ (.A(_05844_),
    .B(_05715_),
    .Y(_05985_));
 sky130_fd_sc_hd__nand3_4 _22628_ (.A(_05983_),
    .B(_05985_),
    .C(_05980_),
    .Y(_05986_));
 sky130_fd_sc_hd__nand2_2 _22629_ (.A(_05861_),
    .B(_05856_),
    .Y(_05987_));
 sky130_fd_sc_hd__a21oi_4 _22630_ (.A1(_05984_),
    .A2(_05986_),
    .B1(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand3_4 _22631_ (.A(_05984_),
    .B(_05986_),
    .C(_05987_),
    .Y(_05989_));
 sky130_fd_sc_hd__and2b_1 _22632_ (.A_N(_05988_),
    .B(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__a21oi_1 _22633_ (.A1(_05868_),
    .A2(_05866_),
    .B1(_05865_),
    .Y(_05991_));
 sky130_fd_sc_hd__xnor2_1 _22634_ (.A(_05990_),
    .B(_05991_),
    .Y(_02636_));
 sky130_fd_sc_hd__nor2_1 _22635_ (.A(_05881_),
    .B(_05888_),
    .Y(_05992_));
 sky130_fd_sc_hd__o21ba_2 _22636_ (.A1(_05877_),
    .A2(_05889_),
    .B1_N(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__nor2_1 _22637_ (.A(_05958_),
    .B(_05964_),
    .Y(_05994_));
 sky130_fd_sc_hd__o21bai_4 _22638_ (.A1(_05953_),
    .A2(_05965_),
    .B1_N(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand3b_1 _22639_ (.A_N(_05885_),
    .B(_05577_),
    .C(_05309_),
    .Y(_05996_));
 sky130_fd_sc_hd__o31a_4 _22640_ (.A1(_14070_),
    .A2(_05418_),
    .A3(_05887_),
    .B1(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__buf_4 _22641_ (.A(_14410_),
    .X(_05998_));
 sky130_fd_sc_hd__nand3b_2 _22642_ (.A_N(_05950_),
    .B(_05361_),
    .C(_05099_),
    .Y(_05999_));
 sky130_fd_sc_hd__o31a_4 _22643_ (.A1(_05878_),
    .A2(_05998_),
    .A3(_05952_),
    .B1(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__clkbuf_4 _22644_ (.A(\pcpi_mul.rs2[6] ),
    .X(_06001_));
 sky130_fd_sc_hd__buf_2 _22645_ (.A(\pcpi_mul.rs1[12] ),
    .X(_06002_));
 sky130_fd_sc_hd__and2_2 _22646_ (.A(_06001_),
    .B(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__nand2_2 _22647_ (.A(_05884_),
    .B(_05320_),
    .Y(_06004_));
 sky130_fd_sc_hd__and2_1 _22648_ (.A(_14061_),
    .B(\pcpi_mul.rs1[10] ),
    .X(_06005_));
 sky130_fd_sc_hd__xor2_4 _22649_ (.A(_06004_),
    .B(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__xor2_4 _22650_ (.A(_06003_),
    .B(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__xnor2_4 _22651_ (.A(_06000_),
    .B(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__xor2_4 _22652_ (.A(_05997_),
    .B(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__xnor2_4 _22653_ (.A(_05995_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__xor2_4 _22654_ (.A(_05993_),
    .B(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__nor2_1 _22655_ (.A(_05893_),
    .B(_05891_),
    .Y(_06012_));
 sky130_fd_sc_hd__a21o_1 _22656_ (.A1(_05873_),
    .A2(_05890_),
    .B1(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__nor2_2 _22657_ (.A(_06011_),
    .B(_06013_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_2 _22658_ (.A(_06013_),
    .B(_06011_),
    .Y(_06015_));
 sky130_vsdinv _22659_ (.A(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__clkbuf_2 _22660_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06017_));
 sky130_fd_sc_hd__clkbuf_4 _22661_ (.A(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__buf_4 _22662_ (.A(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__buf_6 _22663_ (.A(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__nand3b_2 _22664_ (.A_N(_05906_),
    .B(_04879_),
    .C(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__o31ai_4 _22665_ (.A1(_05302_),
    .A2(_14379_),
    .A3(_05908_),
    .B1(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__nor2_1 _22666_ (.A(_05911_),
    .B(_05920_),
    .Y(_06023_));
 sky130_fd_sc_hd__o21bai_4 _22667_ (.A1(_05909_),
    .A2(_05921_),
    .B1_N(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__buf_2 _22668_ (.A(\pcpi_mul.rs2[3] ),
    .X(_06025_));
 sky130_fd_sc_hd__and2_2 _22669_ (.A(_06025_),
    .B(_05770_),
    .X(_06026_));
 sky130_fd_sc_hd__nand2_2 _22670_ (.A(_04904_),
    .B(_06019_),
    .Y(_06027_));
 sky130_fd_sc_hd__buf_2 _22671_ (.A(_14357_),
    .X(_06028_));
 sky130_fd_sc_hd__clkbuf_2 _22672_ (.A(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__buf_2 _22673_ (.A(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__nand2_2 _22674_ (.A(_04876_),
    .B(_06030_),
    .Y(_06031_));
 sky130_fd_sc_hd__xnor2_4 _22675_ (.A(_06027_),
    .B(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__xor2_4 _22676_ (.A(_06026_),
    .B(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__buf_6 _22677_ (.A(_14359_),
    .X(_06034_));
 sky130_fd_sc_hd__nand3b_1 _22678_ (.A_N(_05916_),
    .B(_05117_),
    .C(_05505_),
    .Y(_06035_));
 sky130_fd_sc_hd__o31a_2 _22679_ (.A1(_14097_),
    .A2(_06034_),
    .A3(_05919_),
    .B1(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__clkbuf_4 _22680_ (.A(_14350_),
    .X(_06037_));
 sky130_fd_sc_hd__and2_2 _22681_ (.A(_04713_),
    .B(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__nand2_2 _22682_ (.A(_04924_),
    .B(_05690_),
    .Y(_06039_));
 sky130_fd_sc_hd__buf_2 _22683_ (.A(_14381_),
    .X(_06040_));
 sky130_fd_sc_hd__and2_1 _22684_ (.A(_14073_),
    .B(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__xor2_4 _22685_ (.A(_06039_),
    .B(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__xor2_4 _22686_ (.A(_06038_),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__xnor2_4 _22687_ (.A(_06036_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__xor2_4 _22688_ (.A(_06033_),
    .B(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__xnor2_2 _22689_ (.A(_06024_),
    .B(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__xnor2_2 _22690_ (.A(_06022_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__o21bai_4 _22691_ (.A1(_06014_),
    .A2(_06016_),
    .B1_N(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__nand3b_4 _22692_ (.A_N(_06014_),
    .B(_06047_),
    .C(_06015_),
    .Y(_06049_));
 sky130_fd_sc_hd__nor2_4 _22693_ (.A(_05937_),
    .B(_05967_),
    .Y(_06050_));
 sky130_fd_sc_hd__a21oi_4 _22694_ (.A1(_06048_),
    .A2(_06049_),
    .B1(_06050_),
    .Y(_06051_));
 sky130_vsdinv _22695_ (.A(_06051_),
    .Y(_06052_));
 sky130_fd_sc_hd__nand3_4 _22696_ (.A(_06048_),
    .B(_06050_),
    .C(_06049_),
    .Y(_06053_));
 sky130_fd_sc_hd__a21o_1 _22697_ (.A1(_05892_),
    .A2(_05894_),
    .B1(_05896_),
    .X(_06054_));
 sky130_fd_sc_hd__a21oi_4 _22698_ (.A1(_06054_),
    .A2(_05924_),
    .B1(_05898_),
    .Y(_06055_));
 sky130_vsdinv _22699_ (.A(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__a21o_1 _22700_ (.A1(_06052_),
    .A2(_06053_),
    .B1(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__nand3b_4 _22701_ (.A_N(_06051_),
    .B(_06056_),
    .C(_06053_),
    .Y(_06058_));
 sky130_fd_sc_hd__buf_6 _22702_ (.A(\pcpi_mul.rs2[18] ),
    .X(_06059_));
 sky130_fd_sc_hd__buf_6 _22703_ (.A(_06059_),
    .X(_06060_));
 sky130_fd_sc_hd__buf_4 _22704_ (.A(_06060_),
    .X(_06061_));
 sky130_fd_sc_hd__nand2_4 _22705_ (.A(_06061_),
    .B(_04721_),
    .Y(_06062_));
 sky130_fd_sc_hd__nand2_4 _22706_ (.A(_05966_),
    .B(_05948_),
    .Y(_06063_));
 sky130_fd_sc_hd__or2b_4 _22707_ (.A(_05947_),
    .B_N(_05938_),
    .X(_06064_));
 sky130_fd_sc_hd__o22a_2 _22708_ (.A1(_14454_),
    .A2(_05942_),
    .B1(_05940_),
    .B2(_05946_),
    .X(_06065_));
 sky130_fd_sc_hd__and2_2 _22709_ (.A(_05717_),
    .B(_04974_),
    .X(_06066_));
 sky130_fd_sc_hd__buf_6 _22710_ (.A(_14023_),
    .X(_06067_));
 sky130_fd_sc_hd__nand2_2 _22711_ (.A(_06067_),
    .B(_14448_),
    .Y(_06068_));
 sky130_fd_sc_hd__buf_6 _22712_ (.A(\pcpi_mul.rs2[16] ),
    .X(_06069_));
 sky130_fd_sc_hd__buf_4 _22713_ (.A(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__buf_6 _22714_ (.A(_06070_),
    .X(_06071_));
 sky130_fd_sc_hd__nand2_2 _22715_ (.A(_06071_),
    .B(_04890_),
    .Y(_06072_));
 sky130_fd_sc_hd__xnor2_4 _22716_ (.A(_06068_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__xor2_4 _22717_ (.A(_06066_),
    .B(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__xnor2_4 _22718_ (.A(_06065_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__xor2_4 _22719_ (.A(_06064_),
    .B(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__and2_2 _22720_ (.A(_05355_),
    .B(_05309_),
    .X(_06077_));
 sky130_fd_sc_hd__nand2_2 _22721_ (.A(_14053_),
    .B(_05426_),
    .Y(_06078_));
 sky130_fd_sc_hd__and2_1 _22722_ (.A(_05357_),
    .B(_05046_),
    .X(_06079_));
 sky130_fd_sc_hd__xor2_4 _22723_ (.A(_06078_),
    .B(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__xor2_4 _22724_ (.A(_06077_),
    .B(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__nand3b_2 _22725_ (.A_N(_05961_),
    .B(_14038_),
    .C(_04974_),
    .Y(_06082_));
 sky130_fd_sc_hd__o31a_4 _22726_ (.A1(_14047_),
    .A2(_14428_),
    .A3(_05963_),
    .B1(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__and2_2 _22727_ (.A(_05532_),
    .B(_05091_),
    .X(_06084_));
 sky130_fd_sc_hd__nand2_2 _22728_ (.A(_14041_),
    .B(_05184_),
    .Y(_06085_));
 sky130_fd_sc_hd__and2_1 _22729_ (.A(_05730_),
    .B(_04926_),
    .X(_06086_));
 sky130_fd_sc_hd__xor2_4 _22730_ (.A(_06085_),
    .B(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__xor2_4 _22731_ (.A(_06084_),
    .B(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__xnor2_4 _22732_ (.A(_06083_),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__xnor2_4 _22733_ (.A(_06081_),
    .B(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__xor2_4 _22734_ (.A(_06076_),
    .B(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__xnor2_4 _22735_ (.A(_06063_),
    .B(_06091_),
    .Y(_06092_));
 sky130_fd_sc_hd__xor2_4 _22736_ (.A(_06062_),
    .B(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__nand3_4 _22737_ (.A(_06057_),
    .B(_06058_),
    .C(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__a21oi_2 _22738_ (.A1(_06052_),
    .A2(_06053_),
    .B1(_06056_),
    .Y(_06095_));
 sky130_vsdinv _22739_ (.A(_06058_),
    .Y(_06096_));
 sky130_fd_sc_hd__o21bai_4 _22740_ (.A1(_06095_),
    .A2(_06096_),
    .B1_N(_06093_),
    .Y(_06097_));
 sky130_fd_sc_hd__o2bb2ai_4 _22741_ (.A1_N(_06094_),
    .A2_N(_06097_),
    .B1(_05969_),
    .B2(_05936_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand3b_4 _22742_ (.A_N(_05971_),
    .B(_06097_),
    .C(_06094_),
    .Y(_06099_));
 sky130_fd_sc_hd__and2b_1 _22743_ (.A_N(_05923_),
    .B(_05901_),
    .X(_06100_));
 sky130_fd_sc_hd__a21o_4 _22744_ (.A1(_05922_),
    .A2(_05903_),
    .B1(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__a21o_1 _22745_ (.A1(_05928_),
    .A2(_05933_),
    .B1(_05927_),
    .X(_06102_));
 sky130_fd_sc_hd__xor2_4 _22746_ (.A(_06101_),
    .B(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__a21o_1 _22747_ (.A1(_06098_),
    .A2(_06099_),
    .B1(_06103_),
    .X(_06104_));
 sky130_vsdinv _22748_ (.A(_05974_),
    .Y(_06105_));
 sky130_fd_sc_hd__a21o_1 _22749_ (.A1(_05973_),
    .A2(_05977_),
    .B1(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__nand3_4 _22750_ (.A(_06098_),
    .B(_06103_),
    .C(_06099_),
    .Y(_06107_));
 sky130_fd_sc_hd__nand3_4 _22751_ (.A(_06104_),
    .B(_06106_),
    .C(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__a21oi_2 _22752_ (.A1(_06098_),
    .A2(_06099_),
    .B1(_06103_),
    .Y(_06109_));
 sky130_vsdinv _22753_ (.A(_06107_),
    .Y(_06110_));
 sky130_fd_sc_hd__o21bai_4 _22754_ (.A1(_06109_),
    .A2(_06110_),
    .B1_N(_06106_),
    .Y(_06111_));
 sky130_fd_sc_hd__o2bb2ai_2 _22755_ (.A1_N(_06108_),
    .A2_N(_06111_),
    .B1(_05811_),
    .B2(_05976_),
    .Y(_06112_));
 sky130_fd_sc_hd__nor2_4 _22756_ (.A(_05976_),
    .B(_05811_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand3_4 _22757_ (.A(_06111_),
    .B(_06113_),
    .C(_06108_),
    .Y(_06114_));
 sky130_fd_sc_hd__a21boi_1 _22758_ (.A1(_05983_),
    .A2(_05985_),
    .B1_N(_05980_),
    .Y(_06115_));
 sky130_fd_sc_hd__a21boi_1 _22759_ (.A1(_06112_),
    .A2(_06114_),
    .B1_N(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__nand3b_4 _22760_ (.A_N(_06115_),
    .B(_06114_),
    .C(_06112_),
    .Y(_06117_));
 sky130_fd_sc_hd__and2b_2 _22761_ (.A_N(_06116_),
    .B(_06117_),
    .X(_06118_));
 sky130_vsdinv _22762_ (.A(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__nand3_2 _22763_ (.A(_05862_),
    .B(_05861_),
    .C(_05860_),
    .Y(_06120_));
 sky130_fd_sc_hd__a21oi_4 _22764_ (.A1(_06120_),
    .A2(_05989_),
    .B1(_05988_),
    .Y(_06121_));
 sky130_fd_sc_hd__a31oi_4 _22765_ (.A1(_05868_),
    .A2(_05866_),
    .A3(_05990_),
    .B1(_06121_),
    .Y(_06122_));
 sky130_fd_sc_hd__xor2_1 _22766_ (.A(_06119_),
    .B(_06122_),
    .X(_02637_));
 sky130_fd_sc_hd__nor2_1 _22767_ (.A(_06083_),
    .B(_06088_),
    .Y(_06123_));
 sky130_fd_sc_hd__o21bai_2 _22768_ (.A1(_06081_),
    .A2(_06089_),
    .B1_N(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__nand3b_1 _22769_ (.A_N(_06004_),
    .B(_05577_),
    .C(_05406_),
    .Y(_06125_));
 sky130_fd_sc_hd__o31a_4 _22770_ (.A1(_05576_),
    .A2(_14390_),
    .A3(_06006_),
    .B1(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__buf_4 _22771_ (.A(_14404_),
    .X(_06127_));
 sky130_fd_sc_hd__nand3b_1 _22772_ (.A_N(_06078_),
    .B(_05359_),
    .C(_05101_),
    .Y(_06128_));
 sky130_fd_sc_hd__o31a_4 _22773_ (.A1(_05878_),
    .A2(_06127_),
    .A3(_06080_),
    .B1(_06128_),
    .X(_06129_));
 sky130_fd_sc_hd__and2_2 _22774_ (.A(_06001_),
    .B(_05915_),
    .X(_06130_));
 sky130_fd_sc_hd__nand2_2 _22775_ (.A(_05063_),
    .B(_14387_),
    .Y(_06131_));
 sky130_fd_sc_hd__and2_1 _22776_ (.A(_05130_),
    .B(_05320_),
    .X(_06132_));
 sky130_fd_sc_hd__xor2_4 _22777_ (.A(_06131_),
    .B(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__xor2_4 _22778_ (.A(_06130_),
    .B(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__xnor2_4 _22779_ (.A(_06129_),
    .B(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__xor2_4 _22780_ (.A(_06126_),
    .B(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__xnor2_2 _22781_ (.A(_06124_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__nor2_1 _22782_ (.A(_06000_),
    .B(_06007_),
    .Y(_06138_));
 sky130_fd_sc_hd__o21ba_2 _22783_ (.A1(_05997_),
    .A2(_06008_),
    .B1_N(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__nand2_2 _22784_ (.A(_06137_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__nor2_4 _22785_ (.A(_06139_),
    .B(_06137_),
    .Y(_06141_));
 sky130_vsdinv _22786_ (.A(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__nor2_1 _22787_ (.A(_05993_),
    .B(_06010_),
    .Y(_06143_));
 sky130_fd_sc_hd__a21o_1 _22788_ (.A1(_05995_),
    .A2(_06009_),
    .B1(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__a21o_2 _22789_ (.A1(_06140_),
    .A2(_06142_),
    .B1(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__nand3_4 _22790_ (.A(_06144_),
    .B(_06142_),
    .C(_06140_),
    .Y(_06146_));
 sky130_fd_sc_hd__buf_6 _22791_ (.A(_05913_),
    .X(_06147_));
 sky130_fd_sc_hd__nand3b_2 _22792_ (.A_N(_06027_),
    .B(_05300_),
    .C(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__o31ai_4 _22793_ (.A1(_14088_),
    .A2(_14374_),
    .A3(_06032_),
    .B1(_06148_),
    .Y(_06149_));
 sky130_fd_sc_hd__nor2_1 _22794_ (.A(_06036_),
    .B(_06043_),
    .Y(_06150_));
 sky130_fd_sc_hd__o21bai_4 _22795_ (.A1(_06033_),
    .A2(_06044_),
    .B1_N(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__and2_2 _22796_ (.A(_06025_),
    .B(_06020_),
    .X(_06152_));
 sky130_fd_sc_hd__nand2_2 _22797_ (.A(_04884_),
    .B(_05913_),
    .Y(_06153_));
 sky130_fd_sc_hd__buf_4 _22798_ (.A(_14350_),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_4 _22799_ (.A(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__nand2_2 _22800_ (.A(_04938_),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__xnor2_4 _22801_ (.A(_06153_),
    .B(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__xor2_4 _22802_ (.A(_06152_),
    .B(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__clkbuf_4 _22803_ (.A(_05419_),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_2 _22804_ (.A(_05915_),
    .X(_06160_));
 sky130_fd_sc_hd__buf_4 _22805_ (.A(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__nand3b_1 _22806_ (.A_N(_06039_),
    .B(_06159_),
    .C(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__o31a_2 _22807_ (.A1(_14097_),
    .A2(_14353_),
    .A3(_06042_),
    .B1(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__buf_2 _22808_ (.A(\pcpi_mul.rs1[19] ),
    .X(_06164_));
 sky130_fd_sc_hd__buf_4 _22809_ (.A(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__and2_2 _22810_ (.A(_04713_),
    .B(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__nand2_2 _22811_ (.A(_05109_),
    .B(_05698_),
    .Y(_06167_));
 sky130_fd_sc_hd__and2_1 _22812_ (.A(_04985_),
    .B(_14376_),
    .X(_06168_));
 sky130_fd_sc_hd__xor2_4 _22813_ (.A(_06167_),
    .B(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__xor2_4 _22814_ (.A(_06166_),
    .B(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__xnor2_4 _22815_ (.A(_06163_),
    .B(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__xor2_4 _22816_ (.A(_06158_),
    .B(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__xnor2_4 _22817_ (.A(_06151_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__xnor2_4 _22818_ (.A(_06149_),
    .B(_06173_),
    .Y(_06174_));
 sky130_fd_sc_hd__a21oi_4 _22819_ (.A1(_06145_),
    .A2(_06146_),
    .B1(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__nand3_4 _22820_ (.A(_06145_),
    .B(_06174_),
    .C(_06146_),
    .Y(_06176_));
 sky130_vsdinv _22821_ (.A(_06176_),
    .Y(_06177_));
 sky130_fd_sc_hd__nor2_2 _22822_ (.A(_06063_),
    .B(_06091_),
    .Y(_06178_));
 sky130_fd_sc_hd__o21bai_4 _22823_ (.A1(_06175_),
    .A2(_06177_),
    .B1_N(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__nand3b_4 _22824_ (.A_N(_06175_),
    .B(_06178_),
    .C(_06176_),
    .Y(_06180_));
 sky130_fd_sc_hd__and2_1 _22825_ (.A(_06049_),
    .B(_06015_),
    .X(_06181_));
 sky130_vsdinv _22826_ (.A(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__a21oi_4 _22827_ (.A1(_06179_),
    .A2(_06180_),
    .B1(_06182_),
    .Y(_06183_));
 sky130_fd_sc_hd__nor2_4 _22828_ (.A(_06062_),
    .B(_06092_),
    .Y(_06184_));
 sky130_fd_sc_hd__buf_4 _22829_ (.A(_14013_),
    .X(_06185_));
 sky130_fd_sc_hd__nand2_4 _22830_ (.A(_06185_),
    .B(_04717_),
    .Y(_06186_));
 sky130_fd_sc_hd__nand2_2 _22831_ (.A(_06061_),
    .B(_04874_),
    .Y(_06187_));
 sky130_fd_sc_hd__xnor2_4 _22832_ (.A(_06186_),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__or2_4 _22833_ (.A(_06065_),
    .B(_06074_),
    .X(_06189_));
 sky130_fd_sc_hd__a22o_1 _22834_ (.A1(_05941_),
    .A2(_04969_),
    .B1(_05814_),
    .B2(_04898_),
    .X(_06190_));
 sky130_fd_sc_hd__nand3_4 _22835_ (.A(_05943_),
    .B(_05944_),
    .C(_04890_),
    .Y(_06191_));
 sky130_fd_sc_hd__or2b_1 _22836_ (.A(_06191_),
    .B_N(_04899_),
    .X(_06192_));
 sky130_fd_sc_hd__o2bb2ai_1 _22837_ (.A1_N(_06190_),
    .A2_N(_06192_),
    .B1(_14033_),
    .B2(_14434_),
    .Y(_06193_));
 sky130_fd_sc_hd__o2111ai_4 _22838_ (.A1(_14439_),
    .A2(_06191_),
    .B1(net438),
    .C1(_04929_),
    .D1(_06190_),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_4 _22839_ (.A(_06193_),
    .B(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__o32a_4 _22840_ (.A1(_14033_),
    .A2(_14439_),
    .A3(_06073_),
    .B1(_14445_),
    .B2(_05942_),
    .X(_06196_));
 sky130_fd_sc_hd__xnor2_4 _22841_ (.A(_06195_),
    .B(_06196_),
    .Y(_06197_));
 sky130_fd_sc_hd__xor2_4 _22842_ (.A(_06189_),
    .B(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__and2_2 _22843_ (.A(_05204_),
    .B(_05404_),
    .X(_06199_));
 sky130_fd_sc_hd__buf_6 _22844_ (.A(_05447_),
    .X(_06200_));
 sky130_fd_sc_hd__nand3_4 _22845_ (.A(_05879_),
    .B(_06200_),
    .C(_05106_),
    .Y(_06201_));
 sky130_fd_sc_hd__buf_4 _22846_ (.A(_14053_),
    .X(_06202_));
 sky130_fd_sc_hd__a22o_2 _22847_ (.A1(_05358_),
    .A2(_05427_),
    .B1(_06202_),
    .B2(_05181_),
    .X(_06203_));
 sky130_fd_sc_hd__o21ai_4 _22848_ (.A1(_14405_),
    .A2(_06201_),
    .B1(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__xor2_4 _22849_ (.A(_06199_),
    .B(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__buf_2 _22850_ (.A(_14045_),
    .X(_06206_));
 sky130_fd_sc_hd__buf_4 _22851_ (.A(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__nand3b_1 _22852_ (.A_N(_06085_),
    .B(_05956_),
    .C(_04957_),
    .Y(_06208_));
 sky130_fd_sc_hd__o31a_4 _22853_ (.A1(_06207_),
    .A2(_14422_),
    .A3(_06087_),
    .B1(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__and2_2 _22854_ (.A(_05728_),
    .B(_05429_),
    .X(_06210_));
 sky130_fd_sc_hd__nand2_2 _22855_ (.A(_05732_),
    .B(_05090_),
    .Y(_06211_));
 sky130_fd_sc_hd__and2_2 _22856_ (.A(_05954_),
    .B(_04959_),
    .X(_06212_));
 sky130_fd_sc_hd__xor2_4 _22857_ (.A(_06211_),
    .B(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__xor2_4 _22858_ (.A(_06210_),
    .B(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__xnor2_4 _22859_ (.A(_06209_),
    .B(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__xnor2_4 _22860_ (.A(_06205_),
    .B(_06215_),
    .Y(_06216_));
 sky130_fd_sc_hd__xnor2_4 _22861_ (.A(_06198_),
    .B(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__or2b_1 _22862_ (.A(_06090_),
    .B_N(_06076_),
    .X(_06218_));
 sky130_fd_sc_hd__o21a_2 _22863_ (.A1(_06064_),
    .A2(_06075_),
    .B1(_06218_),
    .X(_06219_));
 sky130_fd_sc_hd__xor2_4 _22864_ (.A(_06217_),
    .B(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__xor2_4 _22865_ (.A(_06188_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__xor2_4 _22866_ (.A(_06184_),
    .B(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__nand3_4 _22867_ (.A(_06182_),
    .B(_06179_),
    .C(_06180_),
    .Y(_06223_));
 sky130_fd_sc_hd__nand3b_4 _22868_ (.A_N(_06183_),
    .B(_06222_),
    .C(_06223_),
    .Y(_06224_));
 sky130_vsdinv _22869_ (.A(_06223_),
    .Y(_06225_));
 sky130_fd_sc_hd__o21bai_4 _22870_ (.A1(_06183_),
    .A2(_06225_),
    .B1_N(_06222_),
    .Y(_06226_));
 sky130_fd_sc_hd__a21bo_1 _22871_ (.A1(_06224_),
    .A2(_06226_),
    .B1_N(_06094_),
    .X(_06227_));
 sky130_fd_sc_hd__nand3b_4 _22872_ (.A_N(_06094_),
    .B(_06226_),
    .C(_06224_),
    .Y(_06228_));
 sky130_fd_sc_hd__or2b_1 _22873_ (.A(_06046_),
    .B_N(_06022_),
    .X(_06229_));
 sky130_fd_sc_hd__a21boi_2 _22874_ (.A1(_06045_),
    .A2(_06024_),
    .B1_N(_06229_),
    .Y(_06230_));
 sky130_vsdinv _22875_ (.A(_06230_),
    .Y(_06231_));
 sky130_fd_sc_hd__o21ai_4 _22876_ (.A1(_06055_),
    .A2(_06051_),
    .B1(_06053_),
    .Y(_06232_));
 sky130_fd_sc_hd__xor2_4 _22877_ (.A(_06231_),
    .B(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__a21oi_2 _22878_ (.A1(_06227_),
    .A2(_06228_),
    .B1(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__nand3_4 _22879_ (.A(_06227_),
    .B(_06233_),
    .C(_06228_),
    .Y(_06235_));
 sky130_vsdinv _22880_ (.A(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__nand2_2 _22881_ (.A(_06107_),
    .B(_06099_),
    .Y(_06237_));
 sky130_fd_sc_hd__o21bai_4 _22882_ (.A1(_06234_),
    .A2(_06236_),
    .B1_N(_06237_),
    .Y(_06238_));
 sky130_fd_sc_hd__a21o_1 _22883_ (.A1(_06227_),
    .A2(_06228_),
    .B1(_06233_),
    .X(_06239_));
 sky130_fd_sc_hd__nand3_4 _22884_ (.A(_06239_),
    .B(_06237_),
    .C(_06235_),
    .Y(_06240_));
 sky130_fd_sc_hd__nand2_1 _22885_ (.A(_06238_),
    .B(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__and2_2 _22886_ (.A(_06102_),
    .B(_06101_),
    .X(_06242_));
 sky130_vsdinv _22887_ (.A(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__nand2_2 _22888_ (.A(_06241_),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__nand3_4 _22889_ (.A(_06238_),
    .B(_06242_),
    .C(_06240_),
    .Y(_06245_));
 sky130_fd_sc_hd__nand2_2 _22890_ (.A(_06114_),
    .B(_06108_),
    .Y(_06246_));
 sky130_fd_sc_hd__a21oi_4 _22891_ (.A1(_06244_),
    .A2(_06245_),
    .B1(_06246_),
    .Y(_06247_));
 sky130_fd_sc_hd__a21boi_2 _22892_ (.A1(_06111_),
    .A2(_06113_),
    .B1_N(_06108_),
    .Y(_06248_));
 sky130_fd_sc_hd__a21oi_2 _22893_ (.A1(_06238_),
    .A2(_06240_),
    .B1(_06242_),
    .Y(_06249_));
 sky130_fd_sc_hd__nor3b_4 _22894_ (.A(_06248_),
    .B(_06249_),
    .C_N(_06245_),
    .Y(_06250_));
 sky130_fd_sc_hd__nor2_8 _22895_ (.A(_06247_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__o21ai_1 _22896_ (.A1(_06119_),
    .A2(_06122_),
    .B1(_06117_),
    .Y(_06252_));
 sky130_fd_sc_hd__xor2_1 _22897_ (.A(_06251_),
    .B(_06252_),
    .X(_02638_));
 sky130_vsdinv _22898_ (.A(_06217_),
    .Y(_06253_));
 sky130_fd_sc_hd__nor2_1 _22899_ (.A(_06219_),
    .B(_06253_),
    .Y(_06254_));
 sky130_vsdinv _22900_ (.A(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__nor2_1 _22901_ (.A(_06129_),
    .B(_06134_),
    .Y(_06256_));
 sky130_fd_sc_hd__o21ba_1 _22902_ (.A1(_06126_),
    .A2(_06135_),
    .B1_N(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__nand3b_1 _22903_ (.A_N(_06131_),
    .B(_05127_),
    .C(_05414_),
    .Y(_06258_));
 sky130_fd_sc_hd__o31a_2 _22904_ (.A1(_14070_),
    .A2(_14384_),
    .A3(_06133_),
    .B1(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__a2bb2oi_4 _22905_ (.A1_N(_06127_),
    .A2_N(_06201_),
    .B1(_06199_),
    .B2(_06203_),
    .Y(_06260_));
 sky130_fd_sc_hd__a22o_1 _22906_ (.A1(_05486_),
    .A2(_05917_),
    .B1(_05063_),
    .B2(_05511_),
    .X(_06261_));
 sky130_fd_sc_hd__nand3_4 _22907_ (.A(_05130_),
    .B(_05162_),
    .C(_14387_),
    .Y(_06262_));
 sky130_fd_sc_hd__or2b_1 _22908_ (.A(_06262_),
    .B_N(_05915_),
    .X(_06263_));
 sky130_fd_sc_hd__buf_4 _22909_ (.A(_14377_),
    .X(_06264_));
 sky130_fd_sc_hd__o2bb2ai_1 _22910_ (.A1_N(_06261_),
    .A2_N(_06263_),
    .B1(_14069_),
    .B2(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__o2111ai_4 _22911_ (.A1(_14382_),
    .A2(_06262_),
    .B1(_04997_),
    .C1(_05610_),
    .D1(_06261_),
    .Y(_06266_));
 sky130_fd_sc_hd__nand2_4 _22912_ (.A(_06265_),
    .B(_06266_),
    .Y(_06267_));
 sky130_fd_sc_hd__xnor2_2 _22913_ (.A(_06260_),
    .B(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__xor2_2 _22914_ (.A(_06259_),
    .B(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__nor2_1 _22915_ (.A(_06209_),
    .B(_06214_),
    .Y(_06270_));
 sky130_fd_sc_hd__o21bai_2 _22916_ (.A1(_06205_),
    .A2(_06215_),
    .B1_N(_06270_),
    .Y(_06271_));
 sky130_fd_sc_hd__xnor2_1 _22917_ (.A(_06269_),
    .B(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__nor2_1 _22918_ (.A(_06257_),
    .B(_06272_),
    .Y(_06273_));
 sky130_vsdinv _22919_ (.A(_06273_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand2_2 _22920_ (.A(_06272_),
    .B(_06257_),
    .Y(_06275_));
 sky130_fd_sc_hd__and2_1 _22921_ (.A(_06136_),
    .B(_06124_),
    .X(_06276_));
 sky130_fd_sc_hd__a211o_2 _22922_ (.A1(_06274_),
    .A2(_06275_),
    .B1(_06276_),
    .C1(_06141_),
    .X(_06277_));
 sky130_fd_sc_hd__o211ai_4 _22923_ (.A1(_06276_),
    .A2(_06141_),
    .B1(_06274_),
    .C1(_06275_),
    .Y(_06278_));
 sky130_fd_sc_hd__buf_2 _22924_ (.A(_06037_),
    .X(_06279_));
 sky130_fd_sc_hd__buf_6 _22925_ (.A(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__nand3b_2 _22926_ (.A_N(_06153_),
    .B(_04947_),
    .C(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__o31ai_4 _22927_ (.A1(_14087_),
    .A2(_14368_),
    .A3(_06157_),
    .B1(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__nor2_1 _22928_ (.A(_06163_),
    .B(_06170_),
    .Y(_06283_));
 sky130_fd_sc_hd__o21bai_4 _22929_ (.A1(_06158_),
    .A2(_06171_),
    .B1_N(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__clkbuf_4 _22930_ (.A(_06029_),
    .X(_06285_));
 sky130_fd_sc_hd__and2_2 _22931_ (.A(_04932_),
    .B(_06285_),
    .X(_06286_));
 sky130_fd_sc_hd__buf_2 _22932_ (.A(_14350_),
    .X(_06287_));
 sky130_fd_sc_hd__buf_4 _22933_ (.A(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__nand2_2 _22934_ (.A(_04904_),
    .B(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__nand2_2 _22935_ (.A(_04909_),
    .B(_06165_),
    .Y(_06290_));
 sky130_fd_sc_hd__xnor2_4 _22936_ (.A(_06289_),
    .B(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__xor2_4 _22937_ (.A(_06286_),
    .B(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__buf_4 _22938_ (.A(_14346_),
    .X(_06293_));
 sky130_fd_sc_hd__nand3b_1 _22939_ (.A_N(_06167_),
    .B(_05117_),
    .C(_05691_),
    .Y(_06294_));
 sky130_fd_sc_hd__o31a_2 _22940_ (.A1(_05056_),
    .A2(_06293_),
    .A3(_06169_),
    .B1(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__clkbuf_4 _22941_ (.A(_14337_),
    .X(_06296_));
 sky130_fd_sc_hd__and2_2 _22942_ (.A(_05045_),
    .B(_06296_),
    .X(_06297_));
 sky130_fd_sc_hd__nand2_2 _22943_ (.A(_05109_),
    .B(_05776_),
    .Y(_06298_));
 sky130_fd_sc_hd__and2_1 _22944_ (.A(_04985_),
    .B(_05698_),
    .X(_06299_));
 sky130_fd_sc_hd__xor2_4 _22945_ (.A(_06298_),
    .B(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__xor2_4 _22946_ (.A(_06297_),
    .B(_06300_),
    .X(_06301_));
 sky130_fd_sc_hd__xnor2_4 _22947_ (.A(_06295_),
    .B(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__xor2_4 _22948_ (.A(_06292_),
    .B(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__xnor2_4 _22949_ (.A(_06284_),
    .B(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__xnor2_4 _22950_ (.A(_06282_),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__a21oi_4 _22951_ (.A1(_06277_),
    .A2(_06278_),
    .B1(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__nand3_4 _22952_ (.A(_06277_),
    .B(_06305_),
    .C(_06278_),
    .Y(_06307_));
 sky130_vsdinv _22953_ (.A(_06307_),
    .Y(_06308_));
 sky130_fd_sc_hd__nor3_4 _22954_ (.A(_06255_),
    .B(_06306_),
    .C(_06308_),
    .Y(_06309_));
 sky130_vsdinv _22955_ (.A(_06309_),
    .Y(_06310_));
 sky130_fd_sc_hd__o21bai_4 _22956_ (.A1(_06306_),
    .A2(_06308_),
    .B1_N(_06254_),
    .Y(_06311_));
 sky130_fd_sc_hd__a21boi_1 _22957_ (.A1(_06145_),
    .A2(_06174_),
    .B1_N(_06146_),
    .Y(_06312_));
 sky130_vsdinv _22958_ (.A(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__a21oi_2 _22959_ (.A1(_06310_),
    .A2(_06311_),
    .B1(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__nand3b_4 _22960_ (.A_N(_06309_),
    .B(_06313_),
    .C(_06311_),
    .Y(_06315_));
 sky130_vsdinv _22961_ (.A(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__nor2_1 _22962_ (.A(_06188_),
    .B(_06220_),
    .Y(_06317_));
 sky130_vsdinv _22963_ (.A(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__buf_2 _22964_ (.A(\pcpi_mul.rs2[18] ),
    .X(_06319_));
 sky130_fd_sc_hd__and2_2 _22965_ (.A(_06319_),
    .B(_04968_),
    .X(_06320_));
 sky130_fd_sc_hd__buf_2 _22966_ (.A(_14008_),
    .X(_06321_));
 sky130_fd_sc_hd__clkbuf_4 _22967_ (.A(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__nand3_4 _22968_ (.A(_06322_),
    .B(_14014_),
    .C(_14448_),
    .Y(_06323_));
 sky130_fd_sc_hd__a22o_2 _22969_ (.A1(_14009_),
    .A2(_04716_),
    .B1(_14014_),
    .B2(_14448_),
    .X(_06324_));
 sky130_fd_sc_hd__o21ai_4 _22970_ (.A1(_14454_),
    .A2(_06323_),
    .B1(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__xnor2_4 _22971_ (.A(_06320_),
    .B(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__or2b_1 _22972_ (.A(_06216_),
    .B_N(_06198_),
    .X(_06327_));
 sky130_fd_sc_hd__o21ai_4 _22973_ (.A1(_06189_),
    .A2(_06197_),
    .B1(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__and2_2 _22974_ (.A(_05354_),
    .B(_05321_),
    .X(_06329_));
 sky130_fd_sc_hd__nand3_4 _22975_ (.A(_05879_),
    .B(_06200_),
    .C(_05516_),
    .Y(_06330_));
 sky130_fd_sc_hd__a22o_2 _22976_ (.A1(_05581_),
    .A2(_05308_),
    .B1(_06202_),
    .B2(_05404_),
    .X(_06331_));
 sky130_fd_sc_hd__o21ai_4 _22977_ (.A1(_05874_),
    .A2(_06330_),
    .B1(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__xnor2_4 _22978_ (.A(_06329_),
    .B(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__a22o_1 _22979_ (.A1(_05634_),
    .A2(_05089_),
    .B1(_05636_),
    .B2(_14414_),
    .X(_06334_));
 sky130_fd_sc_hd__nand3_4 _22980_ (.A(_05954_),
    .B(_14040_),
    .C(_05089_),
    .Y(_06335_));
 sky130_fd_sc_hd__or2b_1 _22981_ (.A(_06335_),
    .B_N(_05586_),
    .X(_06336_));
 sky130_fd_sc_hd__o2bb2ai_2 _22982_ (.A1_N(_06334_),
    .A2_N(_06336_),
    .B1(_14046_),
    .B2(_14410_),
    .Y(_06337_));
 sky130_fd_sc_hd__o2111ai_4 _22983_ (.A1(_14415_),
    .A2(_06335_),
    .B1(_05727_),
    .C1(_05227_),
    .D1(_06334_),
    .Y(_06338_));
 sky130_fd_sc_hd__and2_2 _22984_ (.A(_06337_),
    .B(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__nand3b_1 _22985_ (.A_N(_06211_),
    .B(_05956_),
    .C(_05032_),
    .Y(_06340_));
 sky130_fd_sc_hd__o31a_2 _22986_ (.A1(_06207_),
    .A2(_14417_),
    .A3(_06213_),
    .B1(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__xor2_4 _22987_ (.A(_06339_),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__xor2_4 _22988_ (.A(_06333_),
    .B(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__nor2_4 _22989_ (.A(_06195_),
    .B(_06196_),
    .Y(_06344_));
 sky130_fd_sc_hd__o21a_2 _22990_ (.A1(_14439_),
    .A2(_06191_),
    .B1(_06194_),
    .X(_06345_));
 sky130_fd_sc_hd__buf_4 _22991_ (.A(_06059_),
    .X(_06346_));
 sky130_fd_sc_hd__nand3b_4 _22992_ (.A_N(_06186_),
    .B(_06346_),
    .C(_04908_),
    .Y(_06347_));
 sky130_fd_sc_hd__clkbuf_4 _22993_ (.A(\pcpi_mul.rs2[17] ),
    .X(_06348_));
 sky130_fd_sc_hd__buf_4 _22994_ (.A(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__a22o_2 _22995_ (.A1(_06349_),
    .A2(_05051_),
    .B1(_14027_),
    .B2(_04927_),
    .X(_06350_));
 sky130_fd_sc_hd__clkbuf_4 _22996_ (.A(_06069_),
    .X(_06351_));
 sky130_fd_sc_hd__nand3_4 _22997_ (.A(_06348_),
    .B(_06351_),
    .C(_04897_),
    .Y(_06352_));
 sky130_fd_sc_hd__or2b_1 _22998_ (.A(_06352_),
    .B_N(_04976_),
    .X(_06353_));
 sky130_fd_sc_hd__o2bb2ai_2 _22999_ (.A1_N(_06350_),
    .A2_N(_06353_),
    .B1(_14032_),
    .B2(_14428_),
    .Y(_06354_));
 sky130_fd_sc_hd__buf_4 _23000_ (.A(_05716_),
    .X(_06355_));
 sky130_fd_sc_hd__o2111ai_4 _23001_ (.A1(_05580_),
    .A2(_06352_),
    .B1(_06355_),
    .C1(_05032_),
    .D1(_06350_),
    .Y(_06356_));
 sky130_fd_sc_hd__nand2_2 _23002_ (.A(_06354_),
    .B(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__xnor2_4 _23003_ (.A(_06347_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__xor2_4 _23004_ (.A(_06345_),
    .B(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__xnor2_4 _23005_ (.A(_06344_),
    .B(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__xor2_4 _23006_ (.A(_06343_),
    .B(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__xnor2_4 _23007_ (.A(_06328_),
    .B(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__xor2_4 _23008_ (.A(_06326_),
    .B(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__xor2_4 _23009_ (.A(_06318_),
    .B(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__o21bai_2 _23010_ (.A1(_06314_),
    .A2(_06316_),
    .B1_N(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__nand3b_4 _23011_ (.A_N(_06314_),
    .B(_06364_),
    .C(_06315_),
    .Y(_06366_));
 sky130_fd_sc_hd__and2_1 _23012_ (.A(_06221_),
    .B(_06184_),
    .X(_06367_));
 sky130_vsdinv _23013_ (.A(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__nand2_2 _23014_ (.A(_06224_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__a21o_1 _23015_ (.A1(_06365_),
    .A2(_06366_),
    .B1(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__nand3_4 _23016_ (.A(_06369_),
    .B(_06366_),
    .C(_06365_),
    .Y(_06371_));
 sky130_fd_sc_hd__or2b_1 _23017_ (.A(_06173_),
    .B_N(_06149_),
    .X(_06372_));
 sky130_fd_sc_hd__a21boi_4 _23018_ (.A1(_06172_),
    .A2(_06151_),
    .B1_N(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__a21boi_4 _23019_ (.A1(_06182_),
    .A2(_06179_),
    .B1_N(_06180_),
    .Y(_06374_));
 sky130_fd_sc_hd__xor2_4 _23020_ (.A(_06373_),
    .B(_06374_),
    .X(_06375_));
 sky130_fd_sc_hd__a21oi_1 _23021_ (.A1(_06370_),
    .A2(_06371_),
    .B1(_06375_),
    .Y(_06376_));
 sky130_fd_sc_hd__nand3_4 _23022_ (.A(_06370_),
    .B(_06375_),
    .C(_06371_),
    .Y(_06377_));
 sky130_vsdinv _23023_ (.A(_06377_),
    .Y(_06378_));
 sky130_vsdinv _23024_ (.A(_06233_),
    .Y(_06379_));
 sky130_fd_sc_hd__a21boi_2 _23025_ (.A1(_06226_),
    .A2(_06224_),
    .B1_N(_06094_),
    .Y(_06380_));
 sky130_fd_sc_hd__o21ai_4 _23026_ (.A1(_06379_),
    .A2(_06380_),
    .B1(_06228_),
    .Y(_06381_));
 sky130_fd_sc_hd__o21bai_2 _23027_ (.A1(_06376_),
    .A2(_06378_),
    .B1_N(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2_1 _23028_ (.A(_06370_),
    .B(_06371_),
    .Y(_06383_));
 sky130_vsdinv _23029_ (.A(_06375_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand2_2 _23030_ (.A(_06383_),
    .B(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__nand3_4 _23031_ (.A(_06385_),
    .B(_06381_),
    .C(_06377_),
    .Y(_06386_));
 sky130_fd_sc_hd__and2_1 _23032_ (.A(_06232_),
    .B(_06231_),
    .X(_06387_));
 sky130_fd_sc_hd__a21oi_1 _23033_ (.A1(_06382_),
    .A2(_06386_),
    .B1(_06387_),
    .Y(_06388_));
 sky130_vsdinv _23034_ (.A(_06387_),
    .Y(_06389_));
 sky130_fd_sc_hd__a21oi_4 _23035_ (.A1(_06385_),
    .A2(_06377_),
    .B1(_06381_),
    .Y(_06390_));
 sky130_fd_sc_hd__nor3b_2 _23036_ (.A(_06389_),
    .B(_06390_),
    .C_N(_06386_),
    .Y(_06391_));
 sky130_fd_sc_hd__a21oi_1 _23037_ (.A1(_06239_),
    .A2(_06235_),
    .B1(_06237_),
    .Y(_06392_));
 sky130_fd_sc_hd__o21ai_2 _23038_ (.A1(_06243_),
    .A2(_06392_),
    .B1(_06240_),
    .Y(_06393_));
 sky130_fd_sc_hd__o21bai_1 _23039_ (.A1(_06388_),
    .A2(_06391_),
    .B1_N(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__a21o_1 _23040_ (.A1(_06382_),
    .A2(_06386_),
    .B1(_06387_),
    .X(_06395_));
 sky130_fd_sc_hd__nand3_2 _23041_ (.A(_06382_),
    .B(_06387_),
    .C(_06386_),
    .Y(_06396_));
 sky130_fd_sc_hd__nand3_4 _23042_ (.A(_06395_),
    .B(_06396_),
    .C(_06393_),
    .Y(_06397_));
 sky130_fd_sc_hd__nand2_1 _23043_ (.A(_06394_),
    .B(_06397_),
    .Y(_06398_));
 sky130_vsdinv _23044_ (.A(_05988_),
    .Y(_06399_));
 sky130_fd_sc_hd__nand3_1 _23045_ (.A(_05866_),
    .B(_06399_),
    .C(_05989_),
    .Y(_06400_));
 sky130_fd_sc_hd__nand3b_4 _23046_ (.A_N(_06400_),
    .B(_06118_),
    .C(_06251_),
    .Y(_06401_));
 sky130_vsdinv _23047_ (.A(_06401_),
    .Y(_06402_));
 sky130_fd_sc_hd__nand3_1 _23048_ (.A(_06244_),
    .B(_06246_),
    .C(_06245_),
    .Y(_06403_));
 sky130_fd_sc_hd__o21ai_2 _23049_ (.A1(_06117_),
    .A2(_06247_),
    .B1(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__a31oi_4 _23050_ (.A1(_06118_),
    .A2(_06251_),
    .A3(_06121_),
    .B1(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__a21bo_1 _23051_ (.A1(_05868_),
    .A2(_06402_),
    .B1_N(_06405_),
    .X(_06406_));
 sky130_fd_sc_hd__xnor2_1 _23052_ (.A(_06398_),
    .B(_06406_),
    .Y(_02639_));
 sky130_fd_sc_hd__or2b_1 _23053_ (.A(_06342_),
    .B_N(_06333_),
    .X(_06407_));
 sky130_fd_sc_hd__nand3b_2 _23054_ (.A_N(_06341_),
    .B(_06338_),
    .C(_06337_),
    .Y(_06408_));
 sky130_fd_sc_hd__clkbuf_4 _23055_ (.A(_14384_),
    .X(_06409_));
 sky130_fd_sc_hd__o21a_2 _23056_ (.A1(_06409_),
    .A2(_06262_),
    .B1(_06266_),
    .X(_06410_));
 sky130_fd_sc_hd__a2bb2oi_4 _23057_ (.A1_N(_14400_),
    .A2_N(_06330_),
    .B1(_06329_),
    .B2(_06331_),
    .Y(_06411_));
 sky130_fd_sc_hd__clkbuf_2 _23058_ (.A(\pcpi_mul.rs1[14] ),
    .X(_06412_));
 sky130_fd_sc_hd__a22o_1 _23059_ (.A1(_14062_),
    .A2(_05511_),
    .B1(_14066_),
    .B2(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__nand3_4 _23060_ (.A(_05130_),
    .B(_05162_),
    .C(_14381_),
    .Y(_06414_));
 sky130_fd_sc_hd__or2b_1 _23061_ (.A(_06414_),
    .B_N(_05690_),
    .X(_06415_));
 sky130_fd_sc_hd__o2bb2ai_1 _23062_ (.A1_N(_06413_),
    .A2_N(_06415_),
    .B1(_14069_),
    .B2(_14372_),
    .Y(_06416_));
 sky130_fd_sc_hd__o2111ai_4 _23063_ (.A1(_06264_),
    .A2(_06414_),
    .B1(_04997_),
    .C1(_05699_),
    .D1(_06413_),
    .Y(_06417_));
 sky130_fd_sc_hd__nand2_2 _23064_ (.A(_06416_),
    .B(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__xnor2_1 _23065_ (.A(_06411_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__xor2_1 _23066_ (.A(_06410_),
    .B(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__a21bo_1 _23067_ (.A1(_06407_),
    .A2(_06408_),
    .B1_N(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__nand3b_2 _23068_ (.A_N(_06420_),
    .B(_06408_),
    .C(_06407_),
    .Y(_06422_));
 sky130_fd_sc_hd__nand2_2 _23069_ (.A(_06421_),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__nor2_1 _23070_ (.A(_06260_),
    .B(_06267_),
    .Y(_06424_));
 sky130_fd_sc_hd__o21ba_1 _23071_ (.A1(_06259_),
    .A2(_06268_),
    .B1_N(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__nand2_2 _23072_ (.A(_06423_),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__nor2_1 _23073_ (.A(_06425_),
    .B(_06423_),
    .Y(_06427_));
 sky130_vsdinv _23074_ (.A(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__a21o_1 _23075_ (.A1(_06271_),
    .A2(_06269_),
    .B1(_06273_),
    .X(_06429_));
 sky130_fd_sc_hd__a21o_1 _23076_ (.A1(_06426_),
    .A2(_06428_),
    .B1(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__buf_4 _23077_ (.A(_06164_),
    .X(_06431_));
 sky130_fd_sc_hd__buf_4 _23078_ (.A(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__buf_6 _23079_ (.A(_14085_),
    .X(_06433_));
 sky130_fd_sc_hd__nor3_4 _23080_ (.A(_06433_),
    .B(_14361_),
    .C(_06291_),
    .Y(_06434_));
 sky130_fd_sc_hd__a41oi_4 _23081_ (.A1(_05298_),
    .A2(_05899_),
    .A3(_06432_),
    .A4(_06280_),
    .B1(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__nor2_1 _23082_ (.A(_06295_),
    .B(_06301_),
    .Y(_06436_));
 sky130_fd_sc_hd__o21bai_4 _23083_ (.A1(_06292_),
    .A2(_06302_),
    .B1_N(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__buf_4 _23084_ (.A(_06288_),
    .X(_06438_));
 sky130_fd_sc_hd__and2_2 _23085_ (.A(_06025_),
    .B(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__nand2_2 _23086_ (.A(_04936_),
    .B(_06431_),
    .Y(_06440_));
 sky130_fd_sc_hd__clkbuf_4 _23087_ (.A(_06296_),
    .X(_06441_));
 sky130_fd_sc_hd__nand2_2 _23088_ (.A(_04938_),
    .B(_06441_),
    .Y(_06442_));
 sky130_fd_sc_hd__xnor2_4 _23089_ (.A(_06440_),
    .B(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__xor2_4 _23090_ (.A(_06439_),
    .B(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__clkbuf_4 _23091_ (.A(_04923_),
    .X(_06445_));
 sky130_fd_sc_hd__a22o_1 _23092_ (.A1(_05116_),
    .A2(_06018_),
    .B1(_06445_),
    .B2(_06029_),
    .X(_06446_));
 sky130_fd_sc_hd__nand3_4 _23093_ (.A(_05108_),
    .B(_05050_),
    .C(_05776_),
    .Y(_06447_));
 sky130_fd_sc_hd__or2b_1 _23094_ (.A(_06447_),
    .B_N(_06029_),
    .X(_06448_));
 sky130_fd_sc_hd__o2bb2ai_1 _23095_ (.A1_N(_06446_),
    .A2_N(_06448_),
    .B1(_05056_),
    .B2(_14333_),
    .Y(_06449_));
 sky130_fd_sc_hd__buf_4 _23096_ (.A(_14331_),
    .X(_06450_));
 sky130_fd_sc_hd__o2111ai_4 _23097_ (.A1(_14359_),
    .A2(_06447_),
    .B1(_05319_),
    .C1(_06450_),
    .D1(_06446_),
    .Y(_06451_));
 sky130_fd_sc_hd__and2_2 _23098_ (.A(_06449_),
    .B(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__nand3b_1 _23099_ (.A_N(_06298_),
    .B(_06159_),
    .C(_05700_),
    .Y(_06453_));
 sky130_fd_sc_hd__o31a_2 _23100_ (.A1(_14097_),
    .A2(_14340_),
    .A3(_06300_),
    .B1(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__xor2_4 _23101_ (.A(_06452_),
    .B(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__xor2_4 _23102_ (.A(_06444_),
    .B(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__xnor2_4 _23103_ (.A(_06437_),
    .B(_06456_),
    .Y(_06457_));
 sky130_fd_sc_hd__xor2_4 _23104_ (.A(_06435_),
    .B(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__nand3_4 _23105_ (.A(_06429_),
    .B(_06428_),
    .C(_06426_),
    .Y(_06459_));
 sky130_fd_sc_hd__and3_1 _23106_ (.A(_06430_),
    .B(_06458_),
    .C(_06459_),
    .X(_06460_));
 sky130_vsdinv _23107_ (.A(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__a21o_1 _23108_ (.A1(_06430_),
    .A2(_06459_),
    .B1(_06458_),
    .X(_06462_));
 sky130_fd_sc_hd__and2_1 _23109_ (.A(_06361_),
    .B(_06328_),
    .X(_06463_));
 sky130_fd_sc_hd__a21oi_4 _23110_ (.A1(_06461_),
    .A2(_06462_),
    .B1(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__and3b_2 _23111_ (.A_N(_06460_),
    .B(_06463_),
    .C(_06462_),
    .X(_06465_));
 sky130_fd_sc_hd__o211ai_4 _23112_ (.A1(_06464_),
    .A2(_06465_),
    .B1(_06278_),
    .C1(_06307_),
    .Y(_06466_));
 sky130_fd_sc_hd__a211o_4 _23113_ (.A1(_06278_),
    .A2(_06307_),
    .B1(_06464_),
    .C1(_06465_),
    .X(_06467_));
 sky130_fd_sc_hd__and2b_1 _23114_ (.A_N(_06362_),
    .B(_06326_),
    .X(_06468_));
 sky130_fd_sc_hd__clkbuf_2 _23115_ (.A(\pcpi_mul.rs2[21] ),
    .X(_06469_));
 sky130_fd_sc_hd__buf_4 _23116_ (.A(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__clkbuf_8 _23117_ (.A(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__buf_6 _23118_ (.A(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__and2_2 _23119_ (.A(_06472_),
    .B(_04720_),
    .X(_06473_));
 sky130_fd_sc_hd__and2_2 _23120_ (.A(_06060_),
    .B(_04900_),
    .X(_06474_));
 sky130_fd_sc_hd__nand2_2 _23121_ (.A(_14008_),
    .B(_14447_),
    .Y(_06475_));
 sky130_fd_sc_hd__nand2_2 _23122_ (.A(_14013_),
    .B(_14441_),
    .Y(_06476_));
 sky130_fd_sc_hd__xnor2_4 _23123_ (.A(_06475_),
    .B(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__xor2_4 _23124_ (.A(_06474_),
    .B(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__xor2_4 _23125_ (.A(_06473_),
    .B(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__nand3b_2 _23126_ (.A_N(_06347_),
    .B(_06354_),
    .C(_06356_),
    .Y(_06480_));
 sky130_fd_sc_hd__o21ai_2 _23127_ (.A1(_06345_),
    .A2(_06358_),
    .B1(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__o21a_2 _23128_ (.A1(_14434_),
    .A2(_06352_),
    .B1(_06356_),
    .X(_06482_));
 sky130_fd_sc_hd__a2bb2oi_4 _23129_ (.A1_N(_14452_),
    .A2_N(_06323_),
    .B1(_06320_),
    .B2(_06324_),
    .Y(_06483_));
 sky130_fd_sc_hd__a22o_1 _23130_ (.A1(_06348_),
    .A2(_05111_),
    .B1(_06351_),
    .B2(_05184_),
    .X(_06484_));
 sky130_fd_sc_hd__buf_4 _23131_ (.A(\pcpi_mul.rs2[17] ),
    .X(_06485_));
 sky130_fd_sc_hd__nand3_4 _23132_ (.A(_06485_),
    .B(_06069_),
    .C(_04926_),
    .Y(_06486_));
 sky130_fd_sc_hd__or2b_1 _23133_ (.A(_06486_),
    .B_N(_05959_),
    .X(_06487_));
 sky130_fd_sc_hd__o2bb2ai_1 _23134_ (.A1_N(_06484_),
    .A2_N(_06487_),
    .B1(_14031_),
    .B2(_14422_),
    .Y(_06488_));
 sky130_fd_sc_hd__clkbuf_8 _23135_ (.A(\pcpi_mul.rs2[15] ),
    .X(_06489_));
 sky130_fd_sc_hd__o2111ai_4 _23136_ (.A1(_14427_),
    .A2(_06486_),
    .B1(_06489_),
    .C1(_05091_),
    .D1(_06484_),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_4 _23137_ (.A(_06488_),
    .B(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__xnor2_4 _23138_ (.A(_06483_),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__xor2_4 _23139_ (.A(_06482_),
    .B(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__or2_2 _23140_ (.A(_06481_),
    .B(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__and2_2 _23141_ (.A(_05204_),
    .B(_06002_),
    .X(_06495_));
 sky130_fd_sc_hd__nand3_4 _23142_ (.A(_05358_),
    .B(_05272_),
    .C(_05404_),
    .Y(_06496_));
 sky130_fd_sc_hd__a22o_2 _23143_ (.A1(_05445_),
    .A2(_05613_),
    .B1(_05447_),
    .B2(_05882_),
    .X(_06497_));
 sky130_fd_sc_hd__o21ai_4 _23144_ (.A1(_14393_),
    .A2(_06496_),
    .B1(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__xnor2_4 _23145_ (.A(_06495_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__o21a_2 _23146_ (.A1(_14416_),
    .A2(_06335_),
    .B1(_06338_),
    .X(_06500_));
 sky130_fd_sc_hd__a22o_1 _23147_ (.A1(_14035_),
    .A2(_14414_),
    .B1(_05636_),
    .B2(_14408_),
    .X(_06501_));
 sky130_fd_sc_hd__nand3_4 _23148_ (.A(_14035_),
    .B(\pcpi_mul.rs2[13] ),
    .C(_14414_),
    .Y(_06502_));
 sky130_fd_sc_hd__or2b_1 _23149_ (.A(_06502_),
    .B_N(_05426_),
    .X(_06503_));
 sky130_fd_sc_hd__o2bb2ai_1 _23150_ (.A1_N(_06501_),
    .A2_N(_06503_),
    .B1(_06206_),
    .B2(_14404_),
    .Y(_06504_));
 sky130_fd_sc_hd__o2111ai_4 _23151_ (.A1(_14409_),
    .A2(_06502_),
    .B1(_05727_),
    .C1(_05180_),
    .D1(_06501_),
    .Y(_06505_));
 sky130_fd_sc_hd__nand2_4 _23152_ (.A(_06504_),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__xnor2_2 _23153_ (.A(_06500_),
    .B(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__xnor2_2 _23154_ (.A(_06499_),
    .B(_06507_),
    .Y(_06508_));
 sky130_fd_sc_hd__nand2_2 _23155_ (.A(_06493_),
    .B(_06481_),
    .Y(_06509_));
 sky130_fd_sc_hd__nand3_4 _23156_ (.A(_06494_),
    .B(_06508_),
    .C(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__a21o_1 _23157_ (.A1(_06494_),
    .A2(_06509_),
    .B1(_06508_),
    .X(_06511_));
 sky130_fd_sc_hd__nand2_1 _23158_ (.A(_06359_),
    .B(_06344_),
    .Y(_06512_));
 sky130_fd_sc_hd__o21a_1 _23159_ (.A1(_06343_),
    .A2(_06360_),
    .B1(_06512_),
    .X(_06513_));
 sky130_fd_sc_hd__a21boi_2 _23160_ (.A1(_06510_),
    .A2(_06511_),
    .B1_N(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__and2_1 _23161_ (.A(_06511_),
    .B(_06510_),
    .X(_06515_));
 sky130_fd_sc_hd__nor2b_4 _23162_ (.A(_06513_),
    .B_N(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__nor3_1 _23163_ (.A(_06479_),
    .B(_06514_),
    .C(_06516_),
    .Y(_06517_));
 sky130_vsdinv _23164_ (.A(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__o21ai_2 _23165_ (.A1(_06514_),
    .A2(_06516_),
    .B1(_06479_),
    .Y(_06519_));
 sky130_fd_sc_hd__and3_4 _23166_ (.A(_06468_),
    .B(_06518_),
    .C(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__a21oi_4 _23167_ (.A1(_06518_),
    .A2(_06519_),
    .B1(_06468_),
    .Y(_06521_));
 sky130_fd_sc_hd__o2bb2ai_4 _23168_ (.A1_N(_06466_),
    .A2_N(_06467_),
    .B1(_06520_),
    .B2(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__nor2_4 _23169_ (.A(_06521_),
    .B(_06520_),
    .Y(_06523_));
 sky130_fd_sc_hd__nand3_4 _23170_ (.A(_06467_),
    .B(_06466_),
    .C(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__nor2_1 _23171_ (.A(_06318_),
    .B(_06363_),
    .Y(_06525_));
 sky130_vsdinv _23172_ (.A(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__nand2_2 _23173_ (.A(_06366_),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__a21o_1 _23174_ (.A1(_06522_),
    .A2(_06524_),
    .B1(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__nand3_4 _23175_ (.A(_06527_),
    .B(_06522_),
    .C(_06524_),
    .Y(_06529_));
 sky130_fd_sc_hd__and2b_1 _23176_ (.A_N(_06304_),
    .B(_06282_),
    .X(_06530_));
 sky130_fd_sc_hd__a21o_2 _23177_ (.A1(_06303_),
    .A2(_06284_),
    .B1(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__a21o_1 _23178_ (.A1(_06311_),
    .A2(_06313_),
    .B1(_06309_),
    .X(_06532_));
 sky130_fd_sc_hd__xor2_4 _23179_ (.A(_06531_),
    .B(_06532_),
    .X(_06533_));
 sky130_fd_sc_hd__a21oi_2 _23180_ (.A1(_06528_),
    .A2(_06529_),
    .B1(_06533_),
    .Y(_06534_));
 sky130_vsdinv _23181_ (.A(_06533_),
    .Y(_06535_));
 sky130_fd_sc_hd__a21oi_4 _23182_ (.A1(_06522_),
    .A2(_06524_),
    .B1(_06527_),
    .Y(_06536_));
 sky130_fd_sc_hd__nor3b_4 _23183_ (.A(_06535_),
    .B(_06536_),
    .C_N(_06529_),
    .Y(_06537_));
 sky130_fd_sc_hd__a21oi_1 _23184_ (.A1(_06365_),
    .A2(_06366_),
    .B1(_06369_),
    .Y(_06538_));
 sky130_fd_sc_hd__o21ai_2 _23185_ (.A1(_06384_),
    .A2(_06538_),
    .B1(_06371_),
    .Y(_06539_));
 sky130_fd_sc_hd__o21bai_4 _23186_ (.A1(_06534_),
    .A2(_06537_),
    .B1_N(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__a21o_1 _23187_ (.A1(_06528_),
    .A2(_06529_),
    .B1(_06533_),
    .X(_06541_));
 sky130_fd_sc_hd__nand3_2 _23188_ (.A(_06528_),
    .B(_06533_),
    .C(_06529_),
    .Y(_06542_));
 sky130_fd_sc_hd__nand3_4 _23189_ (.A(_06541_),
    .B(_06542_),
    .C(_06539_),
    .Y(_06543_));
 sky130_fd_sc_hd__a21oi_4 _23190_ (.A1(_06223_),
    .A2(_06180_),
    .B1(_06373_),
    .Y(_06544_));
 sky130_fd_sc_hd__a21oi_1 _23191_ (.A1(_06540_),
    .A2(_06543_),
    .B1(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__nand3_4 _23192_ (.A(_06540_),
    .B(_06544_),
    .C(_06543_),
    .Y(_06546_));
 sky130_vsdinv _23193_ (.A(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__o21ai_4 _23194_ (.A1(_06389_),
    .A2(_06390_),
    .B1(_06386_),
    .Y(_06548_));
 sky130_fd_sc_hd__o21bai_1 _23195_ (.A1(_06545_),
    .A2(_06547_),
    .B1_N(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__o2bb2ai_2 _23196_ (.A1_N(_06543_),
    .A2_N(_06540_),
    .B1(_06374_),
    .B2(_06373_),
    .Y(_06550_));
 sky130_fd_sc_hd__nand3_4 _23197_ (.A(_06550_),
    .B(_06548_),
    .C(_06546_),
    .Y(_06551_));
 sky130_fd_sc_hd__nand2_1 _23198_ (.A(_06549_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__a21boi_1 _23199_ (.A1(_06406_),
    .A2(_06394_),
    .B1_N(_06397_),
    .Y(_06553_));
 sky130_fd_sc_hd__xor2_1 _23200_ (.A(_06552_),
    .B(_06553_),
    .X(_02640_));
 sky130_fd_sc_hd__a31oi_4 _23201_ (.A1(_06467_),
    .A2(_06466_),
    .A3(_06523_),
    .B1(_06520_),
    .Y(_06554_));
 sky130_vsdinv _23202_ (.A(_06516_),
    .Y(_06555_));
 sky130_fd_sc_hd__nor2_1 _23203_ (.A(_06411_),
    .B(_06418_),
    .Y(_06556_));
 sky130_fd_sc_hd__o21ba_1 _23204_ (.A1(_06410_),
    .A2(_06419_),
    .B1_N(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__o21a_2 _23205_ (.A1(_14378_),
    .A2(_06414_),
    .B1(_06417_),
    .X(_06558_));
 sky130_fd_sc_hd__a2bb2oi_4 _23206_ (.A1_N(_14394_),
    .A2_N(_06496_),
    .B1(_06495_),
    .B2(_06497_),
    .Y(_06559_));
 sky130_fd_sc_hd__a22o_1 _23207_ (.A1(_05588_),
    .A2(_14376_),
    .B1(_05884_),
    .B2(_14370_),
    .X(_06560_));
 sky130_fd_sc_hd__nand3_4 _23208_ (.A(_14061_),
    .B(_14065_),
    .C(\pcpi_mul.rs1[14] ),
    .Y(_06561_));
 sky130_fd_sc_hd__or2b_1 _23209_ (.A(_06561_),
    .B_N(_05698_),
    .X(_06562_));
 sky130_fd_sc_hd__o2bb2ai_1 _23210_ (.A1_N(_06560_),
    .A2_N(_06562_),
    .B1(_14069_),
    .B2(_14365_),
    .Y(_06563_));
 sky130_fd_sc_hd__o2111ai_4 _23211_ (.A1(_14371_),
    .A2(_06561_),
    .B1(_06001_),
    .C1(_06018_),
    .D1(_06560_),
    .Y(_06564_));
 sky130_fd_sc_hd__nand2_4 _23212_ (.A(_06563_),
    .B(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__xnor2_2 _23213_ (.A(_06559_),
    .B(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__xor2_2 _23214_ (.A(_06558_),
    .B(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__or2b_1 _23215_ (.A(_06507_),
    .B_N(_06499_),
    .X(_06568_));
 sky130_fd_sc_hd__o21ai_2 _23216_ (.A1(_06506_),
    .A2(_06500_),
    .B1(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__xnor2_1 _23217_ (.A(_06567_),
    .B(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__nor2_1 _23218_ (.A(_06557_),
    .B(_06570_),
    .Y(_06571_));
 sky130_vsdinv _23219_ (.A(_06571_),
    .Y(_06572_));
 sky130_fd_sc_hd__nand2_1 _23220_ (.A(_06570_),
    .B(_06557_),
    .Y(_06573_));
 sky130_fd_sc_hd__o21ai_2 _23221_ (.A1(_06425_),
    .A2(_06423_),
    .B1(_06421_),
    .Y(_06574_));
 sky130_fd_sc_hd__a21o_1 _23222_ (.A1(_06572_),
    .A2(_06573_),
    .B1(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__clkbuf_2 _23223_ (.A(\pcpi_mul.rs1[20] ),
    .X(_06576_));
 sky130_fd_sc_hd__buf_4 _23224_ (.A(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__clkbuf_4 _23225_ (.A(_06577_),
    .X(_06578_));
 sky130_fd_sc_hd__nor3_4 _23226_ (.A(_06433_),
    .B(_14354_),
    .C(_06443_),
    .Y(_06579_));
 sky130_fd_sc_hd__a41oi_4 _23227_ (.A1(_05298_),
    .A2(_05899_),
    .A3(_06578_),
    .A4(_06432_),
    .B1(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__and2b_1 _23228_ (.A_N(_06454_),
    .B(_06452_),
    .X(_06581_));
 sky130_fd_sc_hd__o21bai_4 _23229_ (.A1(_06444_),
    .A2(_06455_),
    .B1_N(_06581_),
    .Y(_06582_));
 sky130_fd_sc_hd__buf_2 _23230_ (.A(_06164_),
    .X(_06583_));
 sky130_fd_sc_hd__buf_4 _23231_ (.A(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__and2_2 _23232_ (.A(_06025_),
    .B(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__nand2_2 _23233_ (.A(_04884_),
    .B(_06577_),
    .Y(_06586_));
 sky130_fd_sc_hd__buf_2 _23234_ (.A(_14331_),
    .X(_06587_));
 sky130_fd_sc_hd__nand2_2 _23235_ (.A(_04876_),
    .B(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__xnor2_4 _23236_ (.A(_06586_),
    .B(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__xor2_4 _23237_ (.A(_06585_),
    .B(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__o21a_2 _23238_ (.A1(_06034_),
    .A2(_06447_),
    .B1(_06451_),
    .X(_06591_));
 sky130_fd_sc_hd__a22o_1 _23239_ (.A1(_05326_),
    .A2(_05912_),
    .B1(_04924_),
    .B2(_06287_),
    .X(_06592_));
 sky130_fd_sc_hd__nand3_4 _23240_ (.A(_05326_),
    .B(_04924_),
    .C(_05912_),
    .Y(_06593_));
 sky130_fd_sc_hd__or2b_1 _23241_ (.A(_06593_),
    .B_N(_06155_),
    .X(_06594_));
 sky130_fd_sc_hd__o2bb2ai_1 _23242_ (.A1_N(_06592_),
    .A2_N(_06594_),
    .B1(_05056_),
    .B2(_14327_),
    .Y(_06595_));
 sky130_fd_sc_hd__buf_4 _23243_ (.A(_14325_),
    .X(_06596_));
 sky130_fd_sc_hd__o2111ai_4 _23244_ (.A1(_14352_),
    .A2(_06593_),
    .B1(_04955_),
    .C1(_06596_),
    .D1(_06592_),
    .Y(_06597_));
 sky130_fd_sc_hd__nand2_4 _23245_ (.A(_06595_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__xnor2_4 _23246_ (.A(_06591_),
    .B(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__xor2_4 _23247_ (.A(_06590_),
    .B(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__xnor2_4 _23248_ (.A(_06582_),
    .B(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__xor2_4 _23249_ (.A(_06580_),
    .B(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__nand3_2 _23250_ (.A(_06572_),
    .B(_06574_),
    .C(_06573_),
    .Y(_06603_));
 sky130_fd_sc_hd__and3_1 _23251_ (.A(_06575_),
    .B(_06602_),
    .C(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__a21o_1 _23252_ (.A1(_06575_),
    .A2(_06603_),
    .B1(_06602_),
    .X(_06605_));
 sky130_fd_sc_hd__nor3b_4 _23253_ (.A(_06555_),
    .B(_06604_),
    .C_N(_06605_),
    .Y(_06606_));
 sky130_vsdinv _23254_ (.A(_06604_),
    .Y(_06607_));
 sky130_fd_sc_hd__a21oi_4 _23255_ (.A1(_06607_),
    .A2(_06605_),
    .B1(_06516_),
    .Y(_06608_));
 sky130_fd_sc_hd__a211o_2 _23256_ (.A1(_06459_),
    .A2(_06461_),
    .B1(_06606_),
    .C1(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__o211ai_4 _23257_ (.A1(_06606_),
    .A2(_06608_),
    .B1(_06459_),
    .C1(_06461_),
    .Y(_06610_));
 sky130_fd_sc_hd__and2_2 _23258_ (.A(_05204_),
    .B(_05511_),
    .X(_06611_));
 sky130_fd_sc_hd__nand3_4 _23259_ (.A(_05445_),
    .B(_05272_),
    .C(_05882_),
    .Y(_06612_));
 sky130_fd_sc_hd__a22o_2 _23260_ (.A1(_14050_),
    .A2(_05882_),
    .B1(_05447_),
    .B2(_05917_),
    .X(_06613_));
 sky130_fd_sc_hd__o21ai_4 _23261_ (.A1(_14388_),
    .A2(_06612_),
    .B1(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__xnor2_4 _23262_ (.A(_06611_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__o21a_2 _23263_ (.A1(_14410_),
    .A2(_06502_),
    .B1(_06505_),
    .X(_06616_));
 sky130_fd_sc_hd__a22o_1 _23264_ (.A1(_05634_),
    .A2(_14408_),
    .B1(_14040_),
    .B2(\pcpi_mul.rs1[9] ),
    .X(_06617_));
 sky130_fd_sc_hd__nand3_4 _23265_ (.A(\pcpi_mul.rs2[14] ),
    .B(\pcpi_mul.rs2[13] ),
    .C(\pcpi_mul.rs1[8] ),
    .Y(_06618_));
 sky130_fd_sc_hd__or2b_1 _23266_ (.A(_06618_),
    .B_N(_05180_),
    .X(_06619_));
 sky130_fd_sc_hd__o2bb2ai_1 _23267_ (.A1_N(_06617_),
    .A2_N(_06619_),
    .B1(_06206_),
    .B2(_14399_),
    .Y(_06620_));
 sky130_fd_sc_hd__o2111ai_4 _23268_ (.A1(_14403_),
    .A2(_06618_),
    .B1(_05727_),
    .C1(_05613_),
    .D1(_06617_),
    .Y(_06621_));
 sky130_fd_sc_hd__nand2_2 _23269_ (.A(_06620_),
    .B(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__xnor2_1 _23270_ (.A(_06616_),
    .B(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__xnor2_1 _23271_ (.A(_06615_),
    .B(_06623_),
    .Y(_06624_));
 sky130_vsdinv _23272_ (.A(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__nor2_1 _23273_ (.A(_06483_),
    .B(_06491_),
    .Y(_06626_));
 sky130_fd_sc_hd__o21bai_4 _23274_ (.A1(_06482_),
    .A2(_06492_),
    .B1_N(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__o21a_2 _23275_ (.A1(_14429_),
    .A2(_06486_),
    .B1(_06490_),
    .X(_06628_));
 sky130_fd_sc_hd__a22o_1 _23276_ (.A1(_14022_),
    .A2(_04959_),
    .B1(_14026_),
    .B2(_14420_),
    .X(_06629_));
 sky130_fd_sc_hd__nand3_4 _23277_ (.A(\pcpi_mul.rs2[17] ),
    .B(_06069_),
    .C(_04959_),
    .Y(_06630_));
 sky130_fd_sc_hd__or2b_1 _23278_ (.A(_06630_),
    .B_N(_05090_),
    .X(_06631_));
 sky130_fd_sc_hd__o2bb2ai_1 _23279_ (.A1_N(_06629_),
    .A2_N(_06631_),
    .B1(_14030_),
    .B2(_14416_),
    .Y(_06632_));
 sky130_fd_sc_hd__o2111ai_4 _23280_ (.A1(_14421_),
    .A2(_06630_),
    .B1(\pcpi_mul.rs2[15] ),
    .C1(_05429_),
    .D1(_06629_),
    .Y(_06633_));
 sky130_fd_sc_hd__and2_2 _23281_ (.A(_06632_),
    .B(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__o32a_4 _23282_ (.A1(_14018_),
    .A2(_14438_),
    .A3(_06477_),
    .B1(_14443_),
    .B2(_06323_),
    .X(_06635_));
 sky130_fd_sc_hd__xor2_4 _23283_ (.A(_06634_),
    .B(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__xor2_4 _23284_ (.A(_06628_),
    .B(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__xnor2_2 _23285_ (.A(_06627_),
    .B(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__nor2_1 _23286_ (.A(_06625_),
    .B(_06638_),
    .Y(_06639_));
 sky130_vsdinv _23287_ (.A(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__nand2_2 _23288_ (.A(_06638_),
    .B(_06625_),
    .Y(_06641_));
 sky130_fd_sc_hd__nand2_2 _23289_ (.A(_06510_),
    .B(_06509_),
    .Y(_06642_));
 sky130_fd_sc_hd__a21oi_4 _23290_ (.A1(_06640_),
    .A2(_06641_),
    .B1(_06642_),
    .Y(_06643_));
 sky130_fd_sc_hd__and3b_2 _23291_ (.A_N(_06639_),
    .B(_06642_),
    .C(_06641_),
    .X(_06644_));
 sky130_fd_sc_hd__nand3b_4 _23292_ (.A_N(_06478_),
    .B(_06472_),
    .C(_04720_),
    .Y(_06645_));
 sky130_fd_sc_hd__clkbuf_4 _23293_ (.A(\pcpi_mul.rs2[22] ),
    .X(_06646_));
 sky130_fd_sc_hd__buf_6 _23294_ (.A(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__nand2_2 _23295_ (.A(_06647_),
    .B(_05533_),
    .Y(_06648_));
 sky130_fd_sc_hd__buf_4 _23296_ (.A(_06469_),
    .X(_06649_));
 sky130_fd_sc_hd__nand2_2 _23297_ (.A(_06649_),
    .B(_04872_),
    .Y(_06650_));
 sky130_fd_sc_hd__xnor2_4 _23298_ (.A(_06648_),
    .B(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__a22o_1 _23299_ (.A1(\pcpi_mul.rs2[20] ),
    .A2(\pcpi_mul.rs1[2] ),
    .B1(\pcpi_mul.rs2[19] ),
    .B2(\pcpi_mul.rs1[3] ),
    .X(_06652_));
 sky130_fd_sc_hd__nand3_4 _23300_ (.A(_14008_),
    .B(\pcpi_mul.rs2[19] ),
    .C(_14441_),
    .Y(_06653_));
 sky130_fd_sc_hd__or2b_1 _23301_ (.A(_06653_),
    .B_N(_04900_),
    .X(_06654_));
 sky130_fd_sc_hd__o2bb2ai_2 _23302_ (.A1_N(_06652_),
    .A2_N(_06654_),
    .B1(_14018_),
    .B2(_14435_),
    .Y(_06655_));
 sky130_fd_sc_hd__o2111ai_4 _23303_ (.A1(_14437_),
    .A2(_06653_),
    .B1(\pcpi_mul.rs2[18] ),
    .C1(_05111_),
    .D1(_06652_),
    .Y(_06656_));
 sky130_fd_sc_hd__nand2_2 _23304_ (.A(_06655_),
    .B(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__xnor2_4 _23305_ (.A(_06651_),
    .B(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__xor2_2 _23306_ (.A(_06645_),
    .B(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__nor3b_4 _23307_ (.A(_06643_),
    .B(_06644_),
    .C_N(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__o21ba_1 _23308_ (.A1(_06643_),
    .A2(_06644_),
    .B1_N(_06659_),
    .X(_06661_));
 sky130_fd_sc_hd__nor3_4 _23309_ (.A(_06518_),
    .B(_06660_),
    .C(_06661_),
    .Y(_06662_));
 sky130_fd_sc_hd__o21a_1 _23310_ (.A1(_06660_),
    .A2(_06661_),
    .B1(_06518_),
    .X(_06663_));
 sky130_fd_sc_hd__nor2_4 _23311_ (.A(_06662_),
    .B(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand3_4 _23312_ (.A(_06609_),
    .B(_06610_),
    .C(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__o2bb2ai_2 _23313_ (.A1_N(_06610_),
    .A2_N(_06609_),
    .B1(_06662_),
    .B2(_06663_),
    .Y(_06666_));
 sky130_fd_sc_hd__nand3b_4 _23314_ (.A_N(_06554_),
    .B(_06665_),
    .C(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__nand2_1 _23315_ (.A(_06666_),
    .B(_06665_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_2 _23316_ (.A(_06554_),
    .B(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__nor2_1 _23317_ (.A(_06435_),
    .B(_06457_),
    .Y(_06670_));
 sky130_fd_sc_hd__a21o_4 _23318_ (.A1(_06456_),
    .A2(_06437_),
    .B1(_06670_),
    .X(_06671_));
 sky130_vsdinv _23319_ (.A(_06465_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand2_2 _23320_ (.A(_06467_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__xor2_4 _23321_ (.A(_06671_),
    .B(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__a21oi_4 _23322_ (.A1(_06667_),
    .A2(_06669_),
    .B1(_06674_),
    .Y(_06675_));
 sky130_fd_sc_hd__nand3_4 _23323_ (.A(_06667_),
    .B(_06674_),
    .C(_06669_),
    .Y(_06676_));
 sky130_vsdinv _23324_ (.A(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__o21ai_2 _23325_ (.A1(_06535_),
    .A2(_06536_),
    .B1(_06529_),
    .Y(_06678_));
 sky130_fd_sc_hd__o21bai_4 _23326_ (.A1(_06675_),
    .A2(_06677_),
    .B1_N(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__nand3b_4 _23327_ (.A_N(_06675_),
    .B(_06676_),
    .C(_06678_),
    .Y(_06680_));
 sky130_fd_sc_hd__a21boi_4 _23328_ (.A1(_06315_),
    .A2(_06310_),
    .B1_N(_06531_),
    .Y(_06681_));
 sky130_fd_sc_hd__a21o_1 _23329_ (.A1(_06679_),
    .A2(_06680_),
    .B1(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__nand3_4 _23330_ (.A(_06679_),
    .B(_06680_),
    .C(_06681_),
    .Y(_06683_));
 sky130_fd_sc_hd__nand2_2 _23331_ (.A(_06546_),
    .B(_06543_),
    .Y(_06684_));
 sky130_fd_sc_hd__a21oi_4 _23332_ (.A1(_06682_),
    .A2(_06683_),
    .B1(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__a21boi_2 _23333_ (.A1(_06540_),
    .A2(_06544_),
    .B1_N(_06543_),
    .Y(_06686_));
 sky130_fd_sc_hd__a21oi_2 _23334_ (.A1(_06679_),
    .A2(_06680_),
    .B1(_06681_),
    .Y(_06687_));
 sky130_fd_sc_hd__nor3b_4 _23335_ (.A(_06686_),
    .B(_06687_),
    .C_N(_06683_),
    .Y(_06688_));
 sky130_fd_sc_hd__nor2_8 _23336_ (.A(_06685_),
    .B(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__nor2_2 _23337_ (.A(_06398_),
    .B(_06552_),
    .Y(_06690_));
 sky130_fd_sc_hd__a21oi_2 _23338_ (.A1(_06550_),
    .A2(_06546_),
    .B1(_06548_),
    .Y(_06691_));
 sky130_fd_sc_hd__a21oi_4 _23339_ (.A1(_06397_),
    .A2(_06551_),
    .B1(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__a21o_1 _23340_ (.A1(_06406_),
    .A2(_06690_),
    .B1(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__xor2_1 _23341_ (.A(_06689_),
    .B(_06693_),
    .X(_02641_));
 sky130_fd_sc_hd__nand2_1 _23342_ (.A(_06637_),
    .B(_06627_),
    .Y(_06694_));
 sky130_fd_sc_hd__o21a_1 _23343_ (.A1(_06625_),
    .A2(_06638_),
    .B1(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__and2_2 _23344_ (.A(_05204_),
    .B(_06412_),
    .X(_06696_));
 sky130_fd_sc_hd__nand3_4 _23345_ (.A(_05358_),
    .B(_06202_),
    .C(_05423_),
    .Y(_06697_));
 sky130_fd_sc_hd__a22o_2 _23346_ (.A1(_05445_),
    .A2(_06002_),
    .B1(_05272_),
    .B2(_06040_),
    .X(_06698_));
 sky130_fd_sc_hd__o21ai_4 _23347_ (.A1(_14383_),
    .A2(_06697_),
    .B1(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__xnor2_4 _23348_ (.A(_06696_),
    .B(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__o21a_2 _23349_ (.A1(_14404_),
    .A2(_06618_),
    .B1(_06621_),
    .X(_06701_));
 sky130_fd_sc_hd__a22o_1 _23350_ (.A1(_05634_),
    .A2(\pcpi_mul.rs1[9] ),
    .B1(_14040_),
    .B2(\pcpi_mul.rs1[10] ),
    .X(_06702_));
 sky130_fd_sc_hd__nand3_4 _23351_ (.A(_14035_),
    .B(_05636_),
    .C(\pcpi_mul.rs1[9] ),
    .Y(_06703_));
 sky130_fd_sc_hd__or2b_1 _23352_ (.A(_06703_),
    .B_N(_14398_),
    .X(_06704_));
 sky130_fd_sc_hd__o2bb2ai_1 _23353_ (.A1_N(_06702_),
    .A2_N(_06704_),
    .B1(_06206_),
    .B2(_14393_),
    .Y(_06705_));
 sky130_fd_sc_hd__o2111ai_4 _23354_ (.A1(_14399_),
    .A2(_06703_),
    .B1(_05440_),
    .C1(_05882_),
    .D1(_06702_),
    .Y(_06706_));
 sky130_fd_sc_hd__nand2_2 _23355_ (.A(_06705_),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__xnor2_1 _23356_ (.A(_06701_),
    .B(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__xnor2_1 _23357_ (.A(_06700_),
    .B(_06708_),
    .Y(_06709_));
 sky130_vsdinv _23358_ (.A(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__o21a_2 _23359_ (.A1(_05057_),
    .A2(_06630_),
    .B1(_06633_),
    .X(_06711_));
 sky130_fd_sc_hd__o21a_2 _23360_ (.A1(_14438_),
    .A2(_06653_),
    .B1(_06656_),
    .X(_06712_));
 sky130_fd_sc_hd__a22o_1 _23361_ (.A1(_14022_),
    .A2(_14420_),
    .B1(_14026_),
    .B2(_05046_),
    .X(_06713_));
 sky130_fd_sc_hd__nand3_4 _23362_ (.A(\pcpi_mul.rs2[17] ),
    .B(_06069_),
    .C(_05089_),
    .Y(_06714_));
 sky130_fd_sc_hd__or2b_1 _23363_ (.A(_06714_),
    .B_N(_05586_),
    .X(_06715_));
 sky130_fd_sc_hd__o2bb2ai_1 _23364_ (.A1_N(_06713_),
    .A2_N(_06715_),
    .B1(_14030_),
    .B2(_14410_),
    .Y(_06716_));
 sky130_fd_sc_hd__o2111ai_4 _23365_ (.A1(_14416_),
    .A2(_06714_),
    .B1(_05716_),
    .C1(_05105_),
    .D1(_06713_),
    .Y(_06717_));
 sky130_fd_sc_hd__nand2_4 _23366_ (.A(_06716_),
    .B(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__xnor2_4 _23367_ (.A(_06712_),
    .B(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__xor2_4 _23368_ (.A(_06711_),
    .B(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__and2b_1 _23369_ (.A_N(_06635_),
    .B(_06634_),
    .X(_06721_));
 sky130_fd_sc_hd__o21bai_2 _23370_ (.A1(_06628_),
    .A2(_06636_),
    .B1_N(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__xnor2_2 _23371_ (.A(_06720_),
    .B(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__nor2_2 _23372_ (.A(_06710_),
    .B(_06723_),
    .Y(_06724_));
 sky130_vsdinv _23373_ (.A(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__nand2_2 _23374_ (.A(_06723_),
    .B(_06710_),
    .Y(_06726_));
 sky130_fd_sc_hd__nor2_4 _23375_ (.A(_06645_),
    .B(_06658_),
    .Y(_06727_));
 sky130_fd_sc_hd__a21oi_4 _23376_ (.A1(_06725_),
    .A2(_06726_),
    .B1(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__nand3b_4 _23377_ (.A_N(_06724_),
    .B(_06727_),
    .C(_06726_),
    .Y(_06729_));
 sky130_fd_sc_hd__nor3b_4 _23378_ (.A(_06695_),
    .B(_06728_),
    .C_N(_06729_),
    .Y(_06730_));
 sky130_vsdinv _23379_ (.A(_06728_),
    .Y(_06731_));
 sky130_vsdinv _23380_ (.A(_06695_),
    .Y(_06732_));
 sky130_fd_sc_hd__a21oi_4 _23381_ (.A1(_06731_),
    .A2(_06729_),
    .B1(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__nand3b_2 _23382_ (.A_N(_06651_),
    .B(_06655_),
    .C(_06656_),
    .Y(_06734_));
 sky130_vsdinv _23383_ (.A(_06734_),
    .Y(_06735_));
 sky130_fd_sc_hd__and2_2 _23384_ (.A(\pcpi_mul.rs2[18] ),
    .B(_04960_),
    .X(_06736_));
 sky130_fd_sc_hd__buf_4 _23385_ (.A(\pcpi_mul.rs2[19] ),
    .X(_06737_));
 sky130_fd_sc_hd__nand3_4 _23386_ (.A(_14009_),
    .B(_06737_),
    .C(_04949_),
    .Y(_06738_));
 sky130_fd_sc_hd__a22o_1 _23387_ (.A1(_06321_),
    .A2(_04897_),
    .B1(_14013_),
    .B2(_05111_),
    .X(_06739_));
 sky130_fd_sc_hd__o21ai_2 _23388_ (.A1(_05580_),
    .A2(_06738_),
    .B1(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__xnor2_2 _23389_ (.A(_06736_),
    .B(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__nand3b_4 _23390_ (.A_N(_06648_),
    .B(_06471_),
    .C(_04908_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_2 _23391_ (.A(_06469_),
    .B(_04890_),
    .Y(_06743_));
 sky130_fd_sc_hd__clkbuf_4 _23392_ (.A(_13997_),
    .X(_06744_));
 sky130_fd_sc_hd__nand3_4 _23393_ (.A(_06744_),
    .B(_14001_),
    .C(_04986_),
    .Y(_06745_));
 sky130_fd_sc_hd__a22o_1 _23394_ (.A1(_13997_),
    .A2(_04716_),
    .B1(_14001_),
    .B2(_04986_),
    .X(_06746_));
 sky130_fd_sc_hd__o21ai_2 _23395_ (.A1(_14452_),
    .A2(_06745_),
    .B1(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__xnor2_2 _23396_ (.A(_06743_),
    .B(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__xnor2_1 _23397_ (.A(_06742_),
    .B(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__xnor2_1 _23398_ (.A(_06741_),
    .B(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__xor2_1 _23399_ (.A(_06735_),
    .B(_06750_),
    .X(_06751_));
 sky130_vsdinv _23400_ (.A(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__o21a_1 _23401_ (.A1(_06730_),
    .A2(_06733_),
    .B1(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__nand3b_1 _23402_ (.A_N(_06728_),
    .B(_06732_),
    .C(_06729_),
    .Y(_06754_));
 sky130_fd_sc_hd__nor3b_4 _23403_ (.A(_06752_),
    .B(_06733_),
    .C_N(_06754_),
    .Y(_06755_));
 sky130_fd_sc_hd__o21ba_1 _23404_ (.A1(_06753_),
    .A2(_06755_),
    .B1_N(_06660_),
    .X(_06756_));
 sky130_vsdinv _23405_ (.A(_06756_),
    .Y(_06757_));
 sky130_vsdinv _23406_ (.A(_06755_),
    .Y(_06758_));
 sky130_fd_sc_hd__nand3b_4 _23407_ (.A_N(_06753_),
    .B(_06758_),
    .C(_06660_),
    .Y(_06759_));
 sky130_fd_sc_hd__buf_4 _23408_ (.A(\pcpi_mul.rs1[21] ),
    .X(_06760_));
 sky130_fd_sc_hd__clkbuf_4 _23409_ (.A(_06760_),
    .X(_06761_));
 sky130_fd_sc_hd__buf_4 _23410_ (.A(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__nor3_4 _23411_ (.A(_14086_),
    .B(_14348_),
    .C(_06589_),
    .Y(_06763_));
 sky130_fd_sc_hd__a41oi_4 _23412_ (.A1(_04946_),
    .A2(_04947_),
    .A3(_06762_),
    .A4(_06578_),
    .B1(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__nor2_1 _23413_ (.A(_06591_),
    .B(_06598_),
    .Y(_06765_));
 sky130_fd_sc_hd__o21bai_4 _23414_ (.A1(_06590_),
    .A2(_06599_),
    .B1_N(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__and2_2 _23415_ (.A(_14082_),
    .B(_06441_),
    .X(_06767_));
 sky130_fd_sc_hd__nand2_2 _23416_ (.A(_04904_),
    .B(_06760_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand2_2 _23417_ (.A(_04909_),
    .B(_06596_),
    .Y(_06769_));
 sky130_fd_sc_hd__xnor2_4 _23418_ (.A(_06768_),
    .B(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__xor2_4 _23419_ (.A(_06767_),
    .B(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__o21a_2 _23420_ (.A1(_14353_),
    .A2(_06593_),
    .B1(_06597_),
    .X(_06772_));
 sky130_fd_sc_hd__a22o_1 _23421_ (.A1(_14073_),
    .A2(_14350_),
    .B1(_05050_),
    .B2(_06164_),
    .X(_06773_));
 sky130_fd_sc_hd__nand3_4 _23422_ (.A(_05108_),
    .B(_05050_),
    .C(_06287_),
    .Y(_06774_));
 sky130_fd_sc_hd__or2b_1 _23423_ (.A(_06774_),
    .B_N(_06583_),
    .X(_06775_));
 sky130_fd_sc_hd__o2bb2ai_1 _23424_ (.A1_N(_06773_),
    .A2_N(_06775_),
    .B1(_14096_),
    .B2(_14320_),
    .Y(_06776_));
 sky130_fd_sc_hd__buf_4 _23425_ (.A(\pcpi_mul.rs1[23] ),
    .X(_06777_));
 sky130_fd_sc_hd__o2111ai_4 _23426_ (.A1(_14345_),
    .A2(_06774_),
    .B1(_05045_),
    .C1(_06777_),
    .D1(_06773_),
    .Y(_06778_));
 sky130_fd_sc_hd__nand2_4 _23427_ (.A(_06776_),
    .B(_06778_),
    .Y(_06779_));
 sky130_fd_sc_hd__xnor2_4 _23428_ (.A(_06772_),
    .B(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__xor2_4 _23429_ (.A(_06771_),
    .B(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__xnor2_4 _23430_ (.A(_06766_),
    .B(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__xor2_4 _23431_ (.A(_06764_),
    .B(_06782_),
    .X(_06783_));
 sky130_vsdinv _23432_ (.A(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__a21o_1 _23433_ (.A1(_06569_),
    .A2(_06567_),
    .B1(_06571_),
    .X(_06785_));
 sky130_fd_sc_hd__o21a_2 _23434_ (.A1(_14372_),
    .A2(_06561_),
    .B1(_06564_),
    .X(_06786_));
 sky130_fd_sc_hd__a2bb2oi_4 _23435_ (.A1_N(_14389_),
    .A2_N(_06612_),
    .B1(_06611_),
    .B2(_06613_),
    .Y(_06787_));
 sky130_fd_sc_hd__a22o_1 _23436_ (.A1(_05130_),
    .A2(_14370_),
    .B1(_05884_),
    .B2(_06017_),
    .X(_06788_));
 sky130_fd_sc_hd__nand3_4 _23437_ (.A(_05129_),
    .B(_14065_),
    .C(\pcpi_mul.rs1[15] ),
    .Y(_06789_));
 sky130_fd_sc_hd__or2b_1 _23438_ (.A(_06789_),
    .B_N(_06017_),
    .X(_06790_));
 sky130_fd_sc_hd__o2bb2ai_1 _23439_ (.A1_N(_06788_),
    .A2_N(_06790_),
    .B1(_14069_),
    .B2(_14358_),
    .Y(_06791_));
 sky130_fd_sc_hd__o2111ai_4 _23440_ (.A1(_14364_),
    .A2(_06789_),
    .B1(_06001_),
    .C1(_05912_),
    .D1(_06788_),
    .Y(_06792_));
 sky130_fd_sc_hd__nand2_4 _23441_ (.A(_06791_),
    .B(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__xnor2_2 _23442_ (.A(_06787_),
    .B(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__xor2_2 _23443_ (.A(_06786_),
    .B(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__or2b_1 _23444_ (.A(_06623_),
    .B_N(_06615_),
    .X(_06796_));
 sky130_fd_sc_hd__o21ai_1 _23445_ (.A1(_06622_),
    .A2(_06616_),
    .B1(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__xnor2_1 _23446_ (.A(_06795_),
    .B(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__nor2_1 _23447_ (.A(_06559_),
    .B(_06565_),
    .Y(_06799_));
 sky130_fd_sc_hd__o21ba_1 _23448_ (.A1(_06558_),
    .A2(_06566_),
    .B1_N(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__nand2_1 _23449_ (.A(_06798_),
    .B(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__nor2_1 _23450_ (.A(_06800_),
    .B(_06798_),
    .Y(_06802_));
 sky130_vsdinv _23451_ (.A(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__and3_2 _23452_ (.A(_06785_),
    .B(_06801_),
    .C(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__a21o_1 _23453_ (.A1(_06801_),
    .A2(_06803_),
    .B1(_06785_),
    .X(_06805_));
 sky130_fd_sc_hd__nor3b_4 _23454_ (.A(_06784_),
    .B(_06804_),
    .C_N(_06805_),
    .Y(_06806_));
 sky130_vsdinv _23455_ (.A(_06806_),
    .Y(_06807_));
 sky130_vsdinv _23456_ (.A(_06804_),
    .Y(_06808_));
 sky130_fd_sc_hd__a21o_1 _23457_ (.A1(_06808_),
    .A2(_06805_),
    .B1(_06783_),
    .X(_06809_));
 sky130_fd_sc_hd__a21oi_4 _23458_ (.A1(_06807_),
    .A2(_06809_),
    .B1(_06644_),
    .Y(_06810_));
 sky130_vsdinv _23459_ (.A(_06644_),
    .Y(_06811_));
 sky130_fd_sc_hd__nor3b_4 _23460_ (.A(_06811_),
    .B(_06806_),
    .C_N(_06809_),
    .Y(_06812_));
 sky130_vsdinv _23461_ (.A(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__a21boi_4 _23462_ (.A1(_06575_),
    .A2(_06602_),
    .B1_N(_06603_),
    .Y(_06814_));
 sky130_vsdinv _23463_ (.A(_06814_),
    .Y(_06815_));
 sky130_fd_sc_hd__nand3b_4 _23464_ (.A_N(_06810_),
    .B(_06813_),
    .C(_06815_),
    .Y(_06816_));
 sky130_fd_sc_hd__o21bai_2 _23465_ (.A1(_06810_),
    .A2(_06812_),
    .B1_N(_06815_),
    .Y(_06817_));
 sky130_fd_sc_hd__a22oi_2 _23466_ (.A1(_06757_),
    .A2(_06759_),
    .B1(_06816_),
    .B2(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__nand2_4 _23467_ (.A(_06757_),
    .B(_06759_),
    .Y(_06819_));
 sky130_fd_sc_hd__nand2_2 _23468_ (.A(_06816_),
    .B(_06817_),
    .Y(_06820_));
 sky130_fd_sc_hd__nor2_4 _23469_ (.A(_06819_),
    .B(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__a31oi_2 _23470_ (.A1(_06609_),
    .A2(_06610_),
    .A3(_06664_),
    .B1(_06662_),
    .Y(_06822_));
 sky130_fd_sc_hd__o21ai_2 _23471_ (.A1(_06818_),
    .A2(_06821_),
    .B1(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__nand3b_2 _23472_ (.A_N(_06819_),
    .B(_06816_),
    .C(_06817_),
    .Y(_06824_));
 sky130_fd_sc_hd__nand2_1 _23473_ (.A(_06820_),
    .B(_06819_),
    .Y(_06825_));
 sky130_fd_sc_hd__nand3b_4 _23474_ (.A_N(_06822_),
    .B(_06824_),
    .C(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__nor2_1 _23475_ (.A(_06580_),
    .B(_06601_),
    .Y(_06827_));
 sky130_fd_sc_hd__a21o_4 _23476_ (.A1(_06600_),
    .A2(_06582_),
    .B1(_06827_),
    .X(_06828_));
 sky130_fd_sc_hd__or2b_2 _23477_ (.A(_06606_),
    .B_N(_06609_),
    .X(_06829_));
 sky130_fd_sc_hd__xor2_4 _23478_ (.A(_06828_),
    .B(_06829_),
    .X(_06830_));
 sky130_fd_sc_hd__a21o_1 _23479_ (.A1(_06823_),
    .A2(_06826_),
    .B1(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__nand3_4 _23480_ (.A(_06823_),
    .B(_06826_),
    .C(_06830_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2_2 _23481_ (.A(_06676_),
    .B(_06667_),
    .Y(_06833_));
 sky130_fd_sc_hd__a21oi_4 _23482_ (.A1(_06831_),
    .A2(_06832_),
    .B1(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__nand3_4 _23483_ (.A(_06833_),
    .B(_06831_),
    .C(_06832_),
    .Y(_06835_));
 sky130_vsdinv _23484_ (.A(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__a21boi_4 _23485_ (.A1(_06467_),
    .A2(_06672_),
    .B1_N(_06671_),
    .Y(_06837_));
 sky130_fd_sc_hd__o21bai_2 _23486_ (.A1(_06834_),
    .A2(_06836_),
    .B1_N(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__nand3b_4 _23487_ (.A_N(_06834_),
    .B(_06837_),
    .C(_06835_),
    .Y(_06839_));
 sky130_fd_sc_hd__nand2_2 _23488_ (.A(_06683_),
    .B(_06680_),
    .Y(_06840_));
 sky130_fd_sc_hd__a21oi_4 _23489_ (.A1(_06838_),
    .A2(_06839_),
    .B1(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__a21boi_2 _23490_ (.A1(_06679_),
    .A2(_06681_),
    .B1_N(_06680_),
    .Y(_06842_));
 sky130_vsdinv _23491_ (.A(_06837_),
    .Y(_06843_));
 sky130_fd_sc_hd__nor3b_4 _23492_ (.A(_06843_),
    .B(_06834_),
    .C_N(_06835_),
    .Y(_06844_));
 sky130_fd_sc_hd__nor3b_4 _23493_ (.A(_06842_),
    .B(_06844_),
    .C_N(_06838_),
    .Y(_06845_));
 sky130_fd_sc_hd__nor2_8 _23494_ (.A(_06841_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__a21oi_1 _23495_ (.A1(_06693_),
    .A2(_06689_),
    .B1(_06688_),
    .Y(_06847_));
 sky130_fd_sc_hd__xnor2_1 _23496_ (.A(_06846_),
    .B(_06847_),
    .Y(_02642_));
 sky130_fd_sc_hd__nor3b_4 _23497_ (.A(_06753_),
    .B(_06755_),
    .C_N(_06660_),
    .Y(_06848_));
 sky130_fd_sc_hd__and2_2 _23498_ (.A(_05204_),
    .B(_05768_),
    .X(_06849_));
 sky130_fd_sc_hd__nand3_4 _23499_ (.A(_05581_),
    .B(_06202_),
    .C(_05512_),
    .Y(_06850_));
 sky130_fd_sc_hd__a22o_2 _23500_ (.A1(_05358_),
    .A2(_06040_),
    .B1(_05272_),
    .B2(_05690_),
    .X(_06851_));
 sky130_fd_sc_hd__o21ai_4 _23501_ (.A1(_06264_),
    .A2(_06850_),
    .B1(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__xnor2_4 _23502_ (.A(_06849_),
    .B(_06852_),
    .Y(_06853_));
 sky130_fd_sc_hd__o21a_2 _23503_ (.A1(_14399_),
    .A2(_06703_),
    .B1(_06706_),
    .X(_06854_));
 sky130_fd_sc_hd__clkbuf_4 _23504_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06855_));
 sky130_fd_sc_hd__a22o_1 _23505_ (.A1(_05954_),
    .A2(\pcpi_mul.rs1[10] ),
    .B1(_06855_),
    .B2(\pcpi_mul.rs1[11] ),
    .X(_06856_));
 sky130_fd_sc_hd__nand3_4 _23506_ (.A(_14035_),
    .B(_05636_),
    .C(\pcpi_mul.rs1[10] ),
    .Y(_06857_));
 sky130_fd_sc_hd__or2b_2 _23507_ (.A(_06857_),
    .B_N(_05320_),
    .X(_06858_));
 sky130_fd_sc_hd__o2bb2ai_1 _23508_ (.A1_N(_06856_),
    .A2_N(_06858_),
    .B1(_06206_),
    .B2(_14388_),
    .Y(_06859_));
 sky130_fd_sc_hd__o2111ai_4 _23509_ (.A1(_14393_),
    .A2(_06857_),
    .B1(_05440_),
    .C1(_05917_),
    .D1(_06856_),
    .Y(_06860_));
 sky130_fd_sc_hd__nand2_2 _23510_ (.A(_06859_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__xnor2_1 _23511_ (.A(_06854_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__xnor2_1 _23512_ (.A(_06853_),
    .B(_06862_),
    .Y(_06863_));
 sky130_vsdinv _23513_ (.A(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__nor2_1 _23514_ (.A(_06712_),
    .B(_06718_),
    .Y(_06865_));
 sky130_fd_sc_hd__o21bai_2 _23515_ (.A1(_06711_),
    .A2(_06719_),
    .B1_N(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__o21a_2 _23516_ (.A1(_05115_),
    .A2(_06714_),
    .B1(_06717_),
    .X(_06867_));
 sky130_fd_sc_hd__a2bb2oi_4 _23517_ (.A1_N(_14433_),
    .A2_N(_06738_),
    .B1(_06736_),
    .B2(_06739_),
    .Y(_06868_));
 sky130_fd_sc_hd__a22o_1 _23518_ (.A1(_14022_),
    .A2(_05046_),
    .B1(_14026_),
    .B2(_05426_),
    .X(_06869_));
 sky130_fd_sc_hd__nand3_4 _23519_ (.A(\pcpi_mul.rs2[17] ),
    .B(_06069_),
    .C(_14414_),
    .Y(_06870_));
 sky130_fd_sc_hd__or2b_1 _23520_ (.A(_06870_),
    .B_N(_05227_),
    .X(_06871_));
 sky130_fd_sc_hd__o2bb2ai_2 _23521_ (.A1_N(_06869_),
    .A2_N(_06871_),
    .B1(_14031_),
    .B2(_14404_),
    .Y(_06872_));
 sky130_fd_sc_hd__o2111ai_4 _23522_ (.A1(_14410_),
    .A2(_06870_),
    .B1(_05716_),
    .C1(_05181_),
    .D1(_06869_),
    .Y(_06873_));
 sky130_fd_sc_hd__nand2_4 _23523_ (.A(_06872_),
    .B(_06873_),
    .Y(_06874_));
 sky130_fd_sc_hd__xnor2_4 _23524_ (.A(_06868_),
    .B(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__xor2_4 _23525_ (.A(_06867_),
    .B(_06875_),
    .X(_06876_));
 sky130_fd_sc_hd__xnor2_2 _23526_ (.A(_06866_),
    .B(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__nor2_2 _23527_ (.A(_06864_),
    .B(_06877_),
    .Y(_06878_));
 sky130_vsdinv _23528_ (.A(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2_2 _23529_ (.A(_06877_),
    .B(_06864_),
    .Y(_06880_));
 sky130_fd_sc_hd__and2_1 _23530_ (.A(_06750_),
    .B(_06735_),
    .X(_06881_));
 sky130_fd_sc_hd__a21o_1 _23531_ (.A1(_06879_),
    .A2(_06880_),
    .B1(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__nand3b_4 _23532_ (.A_N(_06878_),
    .B(_06881_),
    .C(_06880_),
    .Y(_06883_));
 sky130_fd_sc_hd__a21o_1 _23533_ (.A1(_06720_),
    .A2(_06722_),
    .B1(_06724_),
    .X(_06884_));
 sky130_fd_sc_hd__a21oi_4 _23534_ (.A1(_06882_),
    .A2(_06883_),
    .B1(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__and3_1 _23535_ (.A(_06882_),
    .B(_06884_),
    .C(_06883_),
    .X(_06886_));
 sky130_fd_sc_hd__clkbuf_4 _23536_ (.A(\pcpi_mul.rs2[24] ),
    .X(_06887_));
 sky130_fd_sc_hd__buf_4 _23537_ (.A(_06887_),
    .X(_06888_));
 sky130_fd_sc_hd__clkbuf_4 _23538_ (.A(_06888_),
    .X(_06889_));
 sky130_fd_sc_hd__and2_1 _23539_ (.A(_06889_),
    .B(_04720_),
    .X(_06890_));
 sky130_vsdinv _23540_ (.A(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__or2b_1 _23541_ (.A(_06749_),
    .B_N(_06741_),
    .X(_06892_));
 sky130_fd_sc_hd__o21ai_1 _23542_ (.A1(_06742_),
    .A2(_06748_),
    .B1(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__and2_2 _23543_ (.A(_06059_),
    .B(_05099_),
    .X(_06894_));
 sky130_fd_sc_hd__buf_4 _23544_ (.A(_14009_),
    .X(_06895_));
 sky130_fd_sc_hd__buf_4 _23545_ (.A(_14014_),
    .X(_06896_));
 sky130_fd_sc_hd__nand3_4 _23546_ (.A(_06895_),
    .B(_06896_),
    .C(_04928_),
    .Y(_06897_));
 sky130_fd_sc_hd__a22o_2 _23547_ (.A1(_06322_),
    .A2(_04957_),
    .B1(_06185_),
    .B2(_05032_),
    .X(_06898_));
 sky130_fd_sc_hd__o21ai_4 _23548_ (.A1(_05247_),
    .A2(_06897_),
    .B1(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__xor2_4 _23549_ (.A(_06894_),
    .B(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__o22a_2 _23550_ (.A1(_14453_),
    .A2(_06745_),
    .B1(_06743_),
    .B2(_06747_),
    .X(_06901_));
 sky130_fd_sc_hd__and2_2 _23551_ (.A(_06469_),
    .B(_04949_),
    .X(_06902_));
 sky130_fd_sc_hd__nand2_2 _23552_ (.A(_13998_),
    .B(_04906_),
    .Y(_06903_));
 sky130_fd_sc_hd__nand2_2 _23553_ (.A(_06646_),
    .B(_04968_),
    .Y(_06904_));
 sky130_fd_sc_hd__xnor2_4 _23554_ (.A(_06903_),
    .B(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__xor2_4 _23555_ (.A(_06902_),
    .B(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__xnor2_4 _23556_ (.A(_06901_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__xor2_4 _23557_ (.A(_06900_),
    .B(_06907_),
    .X(_06908_));
 sky130_fd_sc_hd__xnor2_1 _23558_ (.A(_06893_),
    .B(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__xor2_1 _23559_ (.A(_06891_),
    .B(_06909_),
    .X(_06910_));
 sky130_vsdinv _23560_ (.A(_06910_),
    .Y(_06911_));
 sky130_fd_sc_hd__o21a_1 _23561_ (.A1(_06885_),
    .A2(_06886_),
    .B1(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__nand3_2 _23562_ (.A(_06882_),
    .B(_06884_),
    .C(_06883_),
    .Y(_06913_));
 sky130_fd_sc_hd__nor3b_4 _23563_ (.A(_06911_),
    .B(_06885_),
    .C_N(_06913_),
    .Y(_06914_));
 sky130_vsdinv _23564_ (.A(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__nand3b_1 _23565_ (.A_N(_06912_),
    .B(_06755_),
    .C(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__o32ai_4 _23566_ (.A1(_06752_),
    .A2(_06730_),
    .A3(_06733_),
    .B1(_06914_),
    .B2(_06912_),
    .Y(_06917_));
 sky130_fd_sc_hd__and2_1 _23567_ (.A(_06916_),
    .B(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__o21a_2 _23568_ (.A1(_14366_),
    .A2(_06789_),
    .B1(_06792_),
    .X(_06919_));
 sky130_fd_sc_hd__a2bb2oi_4 _23569_ (.A1_N(_14383_),
    .A2_N(_06697_),
    .B1(_06696_),
    .B2(_06698_),
    .Y(_06920_));
 sky130_fd_sc_hd__a22o_1 _23570_ (.A1(_05588_),
    .A2(_06017_),
    .B1(_05884_),
    .B2(_14357_),
    .X(_06921_));
 sky130_fd_sc_hd__nand3_4 _23571_ (.A(_14061_),
    .B(_14065_),
    .C(\pcpi_mul.rs1[16] ),
    .Y(_06922_));
 sky130_fd_sc_hd__or2b_1 _23572_ (.A(_06922_),
    .B_N(_06028_),
    .X(_06923_));
 sky130_fd_sc_hd__o2bb2ai_1 _23573_ (.A1_N(_06921_),
    .A2_N(_06923_),
    .B1(_14069_),
    .B2(_14351_),
    .Y(_06924_));
 sky130_fd_sc_hd__o2111ai_4 _23574_ (.A1(_14358_),
    .A2(_06922_),
    .B1(_05483_),
    .C1(_06154_),
    .D1(_06921_),
    .Y(_06925_));
 sky130_fd_sc_hd__nand2_4 _23575_ (.A(_06924_),
    .B(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__xnor2_2 _23576_ (.A(_06920_),
    .B(_06926_),
    .Y(_06927_));
 sky130_fd_sc_hd__xor2_2 _23577_ (.A(_06919_),
    .B(_06927_),
    .X(_06928_));
 sky130_fd_sc_hd__or2b_1 _23578_ (.A(_06708_),
    .B_N(_06700_),
    .X(_06929_));
 sky130_fd_sc_hd__o21ai_2 _23579_ (.A1(_06707_),
    .A2(_06701_),
    .B1(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__xnor2_1 _23580_ (.A(_06928_),
    .B(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__nor2_1 _23581_ (.A(_06787_),
    .B(_06793_),
    .Y(_06932_));
 sky130_fd_sc_hd__o21ba_1 _23582_ (.A1(_06786_),
    .A2(_06794_),
    .B1_N(_06932_),
    .X(_06933_));
 sky130_fd_sc_hd__nand2_2 _23583_ (.A(_06931_),
    .B(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__nor2_1 _23584_ (.A(_06933_),
    .B(_06931_),
    .Y(_06935_));
 sky130_vsdinv _23585_ (.A(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__a21o_1 _23586_ (.A1(_06797_),
    .A2(_06795_),
    .B1(_06802_),
    .X(_06937_));
 sky130_fd_sc_hd__a21o_1 _23587_ (.A1(_06934_),
    .A2(_06936_),
    .B1(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__buf_2 _23588_ (.A(\pcpi_mul.rs1[22] ),
    .X(_06939_));
 sky130_fd_sc_hd__clkbuf_4 _23589_ (.A(_06939_),
    .X(_06940_));
 sky130_fd_sc_hd__buf_4 _23590_ (.A(_06940_),
    .X(_06941_));
 sky130_fd_sc_hd__nor3_4 _23591_ (.A(_14085_),
    .B(_14342_),
    .C(_06770_),
    .Y(_06942_));
 sky130_fd_sc_hd__a41oi_4 _23592_ (.A1(_04886_),
    .A2(_04947_),
    .A3(_06941_),
    .A4(_06762_),
    .B1(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__nor2_1 _23593_ (.A(_06772_),
    .B(_06779_),
    .Y(_06944_));
 sky130_fd_sc_hd__o21bai_4 _23594_ (.A1(_06771_),
    .A2(_06780_),
    .B1_N(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__and2_2 _23595_ (.A(_14082_),
    .B(_06587_),
    .X(_06946_));
 sky130_fd_sc_hd__nand2_2 _23596_ (.A(_14090_),
    .B(_06939_),
    .Y(_06947_));
 sky130_fd_sc_hd__nand2_2 _23597_ (.A(_14093_),
    .B(_06777_),
    .Y(_06948_));
 sky130_fd_sc_hd__xnor2_4 _23598_ (.A(_06947_),
    .B(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__xor2_4 _23599_ (.A(_06946_),
    .B(_06949_),
    .X(_06950_));
 sky130_fd_sc_hd__o21a_2 _23600_ (.A1(_14346_),
    .A2(_06774_),
    .B1(_06778_),
    .X(_06951_));
 sky130_fd_sc_hd__a22o_1 _23601_ (.A1(_05108_),
    .A2(_06164_),
    .B1(_05109_),
    .B2(_06576_),
    .X(_06952_));
 sky130_fd_sc_hd__nand3_4 _23602_ (.A(_04985_),
    .B(_04923_),
    .C(_14344_),
    .Y(_06953_));
 sky130_fd_sc_hd__or2b_2 _23603_ (.A(_06953_),
    .B_N(_06576_),
    .X(_06954_));
 sky130_fd_sc_hd__o2bb2ai_1 _23604_ (.A1_N(_06952_),
    .A2_N(_06954_),
    .B1(_14096_),
    .B2(_14314_),
    .Y(_06955_));
 sky130_fd_sc_hd__clkbuf_2 _23605_ (.A(\pcpi_mul.rs1[24] ),
    .X(_06956_));
 sky130_fd_sc_hd__clkbuf_4 _23606_ (.A(_06956_),
    .X(_06957_));
 sky130_fd_sc_hd__o2111ai_4 _23607_ (.A1(_14338_),
    .A2(_06953_),
    .B1(_04713_),
    .C1(_06957_),
    .D1(_06952_),
    .Y(_06958_));
 sky130_fd_sc_hd__nand2_2 _23608_ (.A(_06955_),
    .B(_06958_),
    .Y(_06959_));
 sky130_fd_sc_hd__xnor2_4 _23609_ (.A(_06951_),
    .B(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__xor2_4 _23610_ (.A(_06950_),
    .B(_06960_),
    .X(_06961_));
 sky130_fd_sc_hd__xnor2_4 _23611_ (.A(_06945_),
    .B(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__xor2_4 _23612_ (.A(_06943_),
    .B(_06962_),
    .X(_06963_));
 sky130_fd_sc_hd__nand3_4 _23613_ (.A(_06937_),
    .B(_06936_),
    .C(_06934_),
    .Y(_06964_));
 sky130_fd_sc_hd__and3_1 _23614_ (.A(_06938_),
    .B(_06963_),
    .C(_06964_),
    .X(_06965_));
 sky130_fd_sc_hd__a21oi_4 _23615_ (.A1(_06938_),
    .A2(_06964_),
    .B1(_06963_),
    .Y(_06966_));
 sky130_vsdinv _23616_ (.A(_06966_),
    .Y(_06967_));
 sky130_fd_sc_hd__o21ai_2 _23617_ (.A1(_06695_),
    .A2(_06728_),
    .B1(_06729_),
    .Y(_06968_));
 sky130_fd_sc_hd__nand3b_4 _23618_ (.A_N(_06965_),
    .B(_06967_),
    .C(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__o21bai_4 _23619_ (.A1(_06966_),
    .A2(_06965_),
    .B1_N(_06968_),
    .Y(_06970_));
 sky130_fd_sc_hd__a21oi_1 _23620_ (.A1(_06805_),
    .A2(_06783_),
    .B1(_06804_),
    .Y(_06971_));
 sky130_vsdinv _23621_ (.A(_06971_),
    .Y(_06972_));
 sky130_fd_sc_hd__a21oi_2 _23622_ (.A1(_06969_),
    .A2(_06970_),
    .B1(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__o211a_1 _23623_ (.A1(_06804_),
    .A2(_06806_),
    .B1(_06970_),
    .C1(_06969_),
    .X(_06974_));
 sky130_fd_sc_hd__nor2_4 _23624_ (.A(_06973_),
    .B(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__nor2_4 _23625_ (.A(_06918_),
    .B(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__and2_1 _23626_ (.A(_06975_),
    .B(_06918_),
    .X(_06977_));
 sky130_fd_sc_hd__nor2_2 _23627_ (.A(_06976_),
    .B(_06977_),
    .Y(_06978_));
 sky130_fd_sc_hd__o21ai_4 _23628_ (.A1(_06848_),
    .A2(_06821_),
    .B1(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__o221ai_4 _23629_ (.A1(_06819_),
    .A2(_06820_),
    .B1(_06976_),
    .B2(_06977_),
    .C1(_06759_),
    .Y(_06980_));
 sky130_fd_sc_hd__nor2_1 _23630_ (.A(_06764_),
    .B(_06782_),
    .Y(_06981_));
 sky130_fd_sc_hd__a21o_4 _23631_ (.A1(_06781_),
    .A2(_06766_),
    .B1(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__o21bai_4 _23632_ (.A1(_06814_),
    .A2(_06810_),
    .B1_N(_06812_),
    .Y(_06983_));
 sky130_fd_sc_hd__xor2_4 _23633_ (.A(_06982_),
    .B(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__a21o_1 _23634_ (.A1(_06979_),
    .A2(_06980_),
    .B1(_06984_),
    .X(_06985_));
 sky130_fd_sc_hd__nand3_4 _23635_ (.A(_06979_),
    .B(_06980_),
    .C(_06984_),
    .Y(_06986_));
 sky130_fd_sc_hd__nand2_2 _23636_ (.A(_06832_),
    .B(_06826_),
    .Y(_06987_));
 sky130_fd_sc_hd__a21o_1 _23637_ (.A1(_06985_),
    .A2(_06986_),
    .B1(_06987_),
    .X(_06988_));
 sky130_fd_sc_hd__nand3_4 _23638_ (.A(_06987_),
    .B(_06985_),
    .C(_06986_),
    .Y(_06989_));
 sky130_fd_sc_hd__and2_2 _23639_ (.A(_06829_),
    .B(_06828_),
    .X(_06990_));
 sky130_fd_sc_hd__a21oi_1 _23640_ (.A1(_06988_),
    .A2(_06989_),
    .B1(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__nand3_4 _23641_ (.A(_06988_),
    .B(_06990_),
    .C(_06989_),
    .Y(_06992_));
 sky130_vsdinv _23642_ (.A(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__o21ai_2 _23643_ (.A1(_06843_),
    .A2(_06834_),
    .B1(_06835_),
    .Y(_06994_));
 sky130_fd_sc_hd__o21bai_1 _23644_ (.A1(_06991_),
    .A2(_06993_),
    .B1_N(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__a21o_1 _23645_ (.A1(_06988_),
    .A2(_06989_),
    .B1(_06990_),
    .X(_06996_));
 sky130_fd_sc_hd__nand3_4 _23646_ (.A(_06996_),
    .B(_06992_),
    .C(_06994_),
    .Y(_06997_));
 sky130_fd_sc_hd__nand2_2 _23647_ (.A(_06995_),
    .B(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__nand3_4 _23648_ (.A(_06690_),
    .B(_06689_),
    .C(_06846_),
    .Y(_06999_));
 sky130_fd_sc_hd__nor2_8 _23649_ (.A(_06999_),
    .B(_06401_),
    .Y(_07000_));
 sky130_fd_sc_hd__nand3_1 _23650_ (.A(_06682_),
    .B(_06684_),
    .C(_06683_),
    .Y(_07001_));
 sky130_fd_sc_hd__nand3_1 _23651_ (.A(_06840_),
    .B(_06838_),
    .C(_06839_),
    .Y(_07002_));
 sky130_fd_sc_hd__o21ai_2 _23652_ (.A1(_07001_),
    .A2(_06841_),
    .B1(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__a31oi_4 _23653_ (.A1(_06846_),
    .A2(_06689_),
    .A3(_06692_),
    .B1(_07003_),
    .Y(_07004_));
 sky130_fd_sc_hd__o21ai_4 _23654_ (.A1(_06999_),
    .A2(_06405_),
    .B1(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__a21oi_4 _23655_ (.A1(_05868_),
    .A2(_07000_),
    .B1(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__xor2_1 _23656_ (.A(_06998_),
    .B(_07006_),
    .X(_02643_));
 sky130_fd_sc_hd__nor2_1 _23657_ (.A(_06920_),
    .B(_06926_),
    .Y(_07007_));
 sky130_fd_sc_hd__o21ba_1 _23658_ (.A1(_06919_),
    .A2(_06927_),
    .B1_N(_07007_),
    .X(_07008_));
 sky130_fd_sc_hd__or2b_1 _23659_ (.A(_06862_),
    .B_N(_06853_),
    .X(_07009_));
 sky130_fd_sc_hd__o21ai_2 _23660_ (.A1(_06861_),
    .A2(_06854_),
    .B1(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__o21a_4 _23661_ (.A1(_06034_),
    .A2(_06922_),
    .B1(_06925_),
    .X(_07011_));
 sky130_fd_sc_hd__a2bb2oi_4 _23662_ (.A1_N(_14378_),
    .A2_N(_06850_),
    .B1(_06849_),
    .B2(_06851_),
    .Y(_07012_));
 sky130_fd_sc_hd__and2_2 _23663_ (.A(_04996_),
    .B(_14344_),
    .X(_07013_));
 sky130_fd_sc_hd__nand2_2 _23664_ (.A(_05162_),
    .B(_14350_),
    .Y(_07014_));
 sky130_fd_sc_hd__and2_1 _23665_ (.A(_05129_),
    .B(\pcpi_mul.rs1[17] ),
    .X(_07015_));
 sky130_fd_sc_hd__xor2_4 _23666_ (.A(_07014_),
    .B(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__xor2_4 _23667_ (.A(_07013_),
    .B(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__xnor2_2 _23668_ (.A(_07012_),
    .B(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__xor2_2 _23669_ (.A(_07011_),
    .B(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__xnor2_1 _23670_ (.A(_07010_),
    .B(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__nor2_1 _23671_ (.A(_07008_),
    .B(_07020_),
    .Y(_07021_));
 sky130_vsdinv _23672_ (.A(_07021_),
    .Y(_07022_));
 sky130_fd_sc_hd__nand2_2 _23673_ (.A(_07020_),
    .B(_07008_),
    .Y(_07023_));
 sky130_fd_sc_hd__a21o_1 _23674_ (.A1(_06930_),
    .A2(_06928_),
    .B1(_06935_),
    .X(_07024_));
 sky130_fd_sc_hd__a21oi_4 _23675_ (.A1(_07022_),
    .A2(_07023_),
    .B1(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__and3_2 _23676_ (.A(_07022_),
    .B(_07024_),
    .C(_07023_),
    .X(_07026_));
 sky130_fd_sc_hd__buf_2 _23677_ (.A(_06777_),
    .X(_07027_));
 sky130_fd_sc_hd__clkbuf_4 _23678_ (.A(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__nor3_4 _23679_ (.A(_06433_),
    .B(_14335_),
    .C(_06949_),
    .Y(_07029_));
 sky130_fd_sc_hd__a41oi_4 _23680_ (.A1(_05298_),
    .A2(_04879_),
    .A3(_07028_),
    .A4(_06941_),
    .B1(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__nor2_1 _23681_ (.A(_06951_),
    .B(_06959_),
    .Y(_07031_));
 sky130_fd_sc_hd__o21bai_4 _23682_ (.A1(_06950_),
    .A2(_06960_),
    .B1_N(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__clkbuf_2 _23683_ (.A(_14325_),
    .X(_07033_));
 sky130_fd_sc_hd__buf_2 _23684_ (.A(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__and2_2 _23685_ (.A(_04932_),
    .B(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__buf_2 _23686_ (.A(_06777_),
    .X(_07036_));
 sky130_fd_sc_hd__nand2_2 _23687_ (.A(_04884_),
    .B(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__clkbuf_4 _23688_ (.A(\pcpi_mul.rs1[24] ),
    .X(_07038_));
 sky130_fd_sc_hd__clkbuf_4 _23689_ (.A(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__nand2_2 _23690_ (.A(_04876_),
    .B(_07039_),
    .Y(_07040_));
 sky130_fd_sc_hd__xnor2_4 _23691_ (.A(_07037_),
    .B(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__xor2_4 _23692_ (.A(_07035_),
    .B(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__nand2_2 _23693_ (.A(_06958_),
    .B(_06954_),
    .Y(_07043_));
 sky130_fd_sc_hd__clkbuf_4 _23694_ (.A(\pcpi_mul.rs1[25] ),
    .X(_07044_));
 sky130_fd_sc_hd__and2_2 _23695_ (.A(_04713_),
    .B(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__buf_6 _23696_ (.A(_14337_),
    .X(_07046_));
 sky130_fd_sc_hd__nand3_4 _23697_ (.A(_05419_),
    .B(_05324_),
    .C(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__buf_2 _23698_ (.A(\pcpi_mul.rs1[21] ),
    .X(_07048_));
 sky130_fd_sc_hd__a22o_2 _23699_ (.A1(_05116_),
    .A2(_06576_),
    .B1(_06445_),
    .B2(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__o21ai_4 _23700_ (.A1(_14332_),
    .A2(_07047_),
    .B1(_07049_),
    .Y(_07050_));
 sky130_fd_sc_hd__xor2_4 _23701_ (.A(_07045_),
    .B(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__xor2_4 _23702_ (.A(_07043_),
    .B(_07051_),
    .X(_07052_));
 sky130_fd_sc_hd__xor2_4 _23703_ (.A(_07042_),
    .B(_07052_),
    .X(_07053_));
 sky130_fd_sc_hd__xnor2_4 _23704_ (.A(_07032_),
    .B(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__xor2_4 _23705_ (.A(_07030_),
    .B(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__nor3b_4 _23706_ (.A(_07025_),
    .B(_07026_),
    .C_N(_07055_),
    .Y(_07056_));
 sky130_vsdinv _23707_ (.A(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__o21bai_2 _23708_ (.A1(_07025_),
    .A2(_07026_),
    .B1_N(_07055_),
    .Y(_07058_));
 sky130_fd_sc_hd__nand2_2 _23709_ (.A(_06913_),
    .B(_06883_),
    .Y(_07059_));
 sky130_fd_sc_hd__a21o_1 _23710_ (.A1(_07057_),
    .A2(_07058_),
    .B1(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__nand3b_4 _23711_ (.A_N(_07056_),
    .B(_07059_),
    .C(_07058_),
    .Y(_07061_));
 sky130_fd_sc_hd__a21boi_2 _23712_ (.A1(_06938_),
    .A2(_06963_),
    .B1_N(_06964_),
    .Y(_07062_));
 sky130_fd_sc_hd__a21bo_1 _23713_ (.A1(_07060_),
    .A2(_07061_),
    .B1_N(_07062_),
    .X(_07063_));
 sky130_fd_sc_hd__nand3b_4 _23714_ (.A_N(_07062_),
    .B(_07060_),
    .C(_07061_),
    .Y(_07064_));
 sky130_fd_sc_hd__and2_2 _23715_ (.A(_05205_),
    .B(_05777_),
    .X(_07065_));
 sky130_fd_sc_hd__nand2_2 _23716_ (.A(_05271_),
    .B(_14370_),
    .Y(_07066_));
 sky130_fd_sc_hd__and2_1 _23717_ (.A(\pcpi_mul.rs2[11] ),
    .B(\pcpi_mul.rs1[14] ),
    .X(_07067_));
 sky130_fd_sc_hd__xor2_4 _23718_ (.A(_07066_),
    .B(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__xnor2_4 _23719_ (.A(_07065_),
    .B(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__nand2_2 _23720_ (.A(_06860_),
    .B(_06858_),
    .Y(_07070_));
 sky130_fd_sc_hd__and2_2 _23721_ (.A(_05727_),
    .B(_05511_),
    .X(_07071_));
 sky130_fd_sc_hd__nand2_2 _23722_ (.A(_14040_),
    .B(\pcpi_mul.rs1[12] ),
    .Y(_07072_));
 sky130_fd_sc_hd__and2_1 _23723_ (.A(\pcpi_mul.rs2[14] ),
    .B(\pcpi_mul.rs1[11] ),
    .X(_07073_));
 sky130_fd_sc_hd__xor2_4 _23724_ (.A(_07072_),
    .B(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__xor2_4 _23725_ (.A(_07071_),
    .B(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__xor2_4 _23726_ (.A(_07070_),
    .B(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__xnor2_2 _23727_ (.A(_07069_),
    .B(_07076_),
    .Y(_07077_));
 sky130_vsdinv _23728_ (.A(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__nor2_1 _23729_ (.A(_06868_),
    .B(_06874_),
    .Y(_07079_));
 sky130_fd_sc_hd__o21bai_2 _23730_ (.A1(_06867_),
    .A2(_06875_),
    .B1_N(_07079_),
    .Y(_07080_));
 sky130_fd_sc_hd__o21a_2 _23731_ (.A1(_14412_),
    .A2(_06870_),
    .B1(_06873_),
    .X(_07081_));
 sky130_fd_sc_hd__a2bb2oi_4 _23732_ (.A1_N(_05247_),
    .A2_N(_06897_),
    .B1(_06894_),
    .B2(_06898_),
    .Y(_07082_));
 sky130_fd_sc_hd__and2_2 _23733_ (.A(_06489_),
    .B(_05241_),
    .X(_07083_));
 sky130_fd_sc_hd__nand2_2 _23734_ (.A(_06351_),
    .B(_05236_),
    .Y(_07084_));
 sky130_fd_sc_hd__and2_1 _23735_ (.A(_06485_),
    .B(_05426_),
    .X(_07085_));
 sky130_fd_sc_hd__xor2_4 _23736_ (.A(_07084_),
    .B(_07085_),
    .X(_07086_));
 sky130_fd_sc_hd__xor2_4 _23737_ (.A(_07083_),
    .B(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__xnor2_2 _23738_ (.A(_07082_),
    .B(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__xor2_2 _23739_ (.A(_07081_),
    .B(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__xnor2_1 _23740_ (.A(_07080_),
    .B(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__nor2_1 _23741_ (.A(_07078_),
    .B(_07090_),
    .Y(_07091_));
 sky130_fd_sc_hd__and2_1 _23742_ (.A(_06908_),
    .B(_06893_),
    .X(_07092_));
 sky130_fd_sc_hd__nand2_1 _23743_ (.A(_07090_),
    .B(_07078_),
    .Y(_07093_));
 sky130_fd_sc_hd__and3b_1 _23744_ (.A_N(_07091_),
    .B(_07092_),
    .C(_07093_),
    .X(_07094_));
 sky130_vsdinv _23745_ (.A(_07094_),
    .Y(_07095_));
 sky130_vsdinv _23746_ (.A(_07091_),
    .Y(_07096_));
 sky130_fd_sc_hd__a21o_1 _23747_ (.A1(_07096_),
    .A2(_07093_),
    .B1(_07092_),
    .X(_07097_));
 sky130_fd_sc_hd__a21o_1 _23748_ (.A1(_06876_),
    .A2(_06866_),
    .B1(_06878_),
    .X(_07098_));
 sky130_fd_sc_hd__a21o_1 _23749_ (.A1(_07095_),
    .A2(_07097_),
    .B1(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__nand3b_4 _23750_ (.A_N(_07094_),
    .B(_07098_),
    .C(_07097_),
    .Y(_07100_));
 sky130_fd_sc_hd__buf_2 _23751_ (.A(\pcpi_mul.rs2[25] ),
    .X(_07101_));
 sky130_fd_sc_hd__buf_4 _23752_ (.A(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__buf_4 _23753_ (.A(_07102_),
    .X(_07103_));
 sky130_fd_sc_hd__buf_8 _23754_ (.A(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__nand2_4 _23755_ (.A(_07104_),
    .B(_04718_),
    .Y(_07105_));
 sky130_fd_sc_hd__buf_4 _23756_ (.A(\pcpi_mul.rs2[24] ),
    .X(_07106_));
 sky130_fd_sc_hd__buf_6 _23757_ (.A(_07106_),
    .X(_07107_));
 sky130_fd_sc_hd__nand2_1 _23758_ (.A(_07107_),
    .B(_04873_),
    .Y(_07108_));
 sky130_fd_sc_hd__xor2_1 _23759_ (.A(_07105_),
    .B(_07108_),
    .X(_07109_));
 sky130_vsdinv _23760_ (.A(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__nor2_1 _23761_ (.A(_06901_),
    .B(_06906_),
    .Y(_07111_));
 sky130_fd_sc_hd__o21bai_4 _23762_ (.A1(_06900_),
    .A2(_06907_),
    .B1_N(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__and2_2 _23763_ (.A(_06346_),
    .B(_05191_),
    .X(_07113_));
 sky130_fd_sc_hd__nand2_2 _23764_ (.A(_14013_),
    .B(_05090_),
    .Y(_07114_));
 sky130_fd_sc_hd__and2_1 _23765_ (.A(_14008_),
    .B(_14426_),
    .X(_07115_));
 sky130_fd_sc_hd__xor2_4 _23766_ (.A(_07114_),
    .B(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__xor2_4 _23767_ (.A(_07113_),
    .B(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__and2_2 _23768_ (.A(_06469_),
    .B(_04976_),
    .X(_07118_));
 sky130_fd_sc_hd__nand2_2 _23769_ (.A(_06646_),
    .B(_05051_),
    .Y(_07119_));
 sky130_fd_sc_hd__and2_2 _23770_ (.A(_06744_),
    .B(_04988_),
    .X(_07120_));
 sky130_fd_sc_hd__xor2_4 _23771_ (.A(_07119_),
    .B(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__xor2_4 _23772_ (.A(_07118_),
    .B(_07121_),
    .X(_07122_));
 sky130_fd_sc_hd__clkbuf_4 _23773_ (.A(_14004_),
    .X(_07123_));
 sky130_fd_sc_hd__o32a_4 _23774_ (.A1(_07123_),
    .A2(_05178_),
    .A3(_06905_),
    .B1(_14444_),
    .B2(_06745_),
    .X(_07124_));
 sky130_fd_sc_hd__xnor2_4 _23775_ (.A(_07122_),
    .B(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__xor2_4 _23776_ (.A(_07117_),
    .B(_07125_),
    .X(_07126_));
 sky130_fd_sc_hd__xnor2_4 _23777_ (.A(_07112_),
    .B(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__nor2_8 _23778_ (.A(_07110_),
    .B(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__and2_1 _23779_ (.A(_07127_),
    .B(_07110_),
    .X(_07129_));
 sky130_fd_sc_hd__nor2_1 _23780_ (.A(_06891_),
    .B(_06909_),
    .Y(_07130_));
 sky130_fd_sc_hd__nor3b_4 _23781_ (.A(_07128_),
    .B(_07129_),
    .C_N(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__o21ba_1 _23782_ (.A1(_07128_),
    .A2(_07129_),
    .B1_N(_07130_),
    .X(_07132_));
 sky130_fd_sc_hd__nor2_4 _23783_ (.A(_07131_),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__a21oi_4 _23784_ (.A1(_07099_),
    .A2(_07100_),
    .B1(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__nand3_1 _23785_ (.A(_07099_),
    .B(_07133_),
    .C(_07100_),
    .Y(_07135_));
 sky130_vsdinv _23786_ (.A(_07135_),
    .Y(_07136_));
 sky130_fd_sc_hd__nor3_4 _23787_ (.A(_06915_),
    .B(_07134_),
    .C(_07136_),
    .Y(_07137_));
 sky130_vsdinv _23788_ (.A(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__o21bai_4 _23789_ (.A1(_07134_),
    .A2(_07136_),
    .B1_N(_06914_),
    .Y(_07139_));
 sky130_fd_sc_hd__a22oi_2 _23790_ (.A1(_07063_),
    .A2(_07064_),
    .B1(_07138_),
    .B2(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__nand2_1 _23791_ (.A(_07063_),
    .B(_07064_),
    .Y(_07141_));
 sky130_fd_sc_hd__nand2_1 _23792_ (.A(_07138_),
    .B(_07139_),
    .Y(_07142_));
 sky130_fd_sc_hd__nor2_1 _23793_ (.A(_07141_),
    .B(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__a21boi_1 _23794_ (.A1(_06975_),
    .A2(_06917_),
    .B1_N(_06916_),
    .Y(_07144_));
 sky130_vsdinv _23795_ (.A(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__o21bai_2 _23796_ (.A1(_07140_),
    .A2(_07143_),
    .B1_N(_07145_),
    .Y(_07146_));
 sky130_fd_sc_hd__nand3b_2 _23797_ (.A_N(_07141_),
    .B(_07138_),
    .C(_07139_),
    .Y(_07147_));
 sky130_fd_sc_hd__nand2_1 _23798_ (.A(_07142_),
    .B(_07141_),
    .Y(_07148_));
 sky130_fd_sc_hd__nand3_4 _23799_ (.A(_07147_),
    .B(_07148_),
    .C(_07145_),
    .Y(_07149_));
 sky130_fd_sc_hd__nand2_1 _23800_ (.A(_07146_),
    .B(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__nor2_2 _23801_ (.A(_06943_),
    .B(_06962_),
    .Y(_07151_));
 sky130_fd_sc_hd__a21oi_4 _23802_ (.A1(_06961_),
    .A2(_06945_),
    .B1(_07151_),
    .Y(_07152_));
 sky130_fd_sc_hd__a21boi_4 _23803_ (.A1(_06972_),
    .A2(_06970_),
    .B1_N(_06969_),
    .Y(_07153_));
 sky130_fd_sc_hd__xor2_4 _23804_ (.A(_07152_),
    .B(_07153_),
    .X(_07154_));
 sky130_vsdinv _23805_ (.A(_07154_),
    .Y(_07155_));
 sky130_fd_sc_hd__nand2_2 _23806_ (.A(_07150_),
    .B(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__nand3_4 _23807_ (.A(_07146_),
    .B(_07149_),
    .C(_07154_),
    .Y(_07157_));
 sky130_fd_sc_hd__nand2_2 _23808_ (.A(_06986_),
    .B(_06979_),
    .Y(_07158_));
 sky130_fd_sc_hd__a21oi_2 _23809_ (.A1(_07156_),
    .A2(_07157_),
    .B1(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__nand3_4 _23810_ (.A(_07156_),
    .B(_07158_),
    .C(_07157_),
    .Y(_07160_));
 sky130_vsdinv _23811_ (.A(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__and2_1 _23812_ (.A(_06983_),
    .B(_06982_),
    .X(_07162_));
 sky130_fd_sc_hd__o21bai_2 _23813_ (.A1(_07159_),
    .A2(_07161_),
    .B1_N(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__nand3b_4 _23814_ (.A_N(_07159_),
    .B(_07162_),
    .C(_07160_),
    .Y(_07164_));
 sky130_fd_sc_hd__nand2_1 _23815_ (.A(_07163_),
    .B(_07164_),
    .Y(_07165_));
 sky130_vsdinv _23816_ (.A(_06990_),
    .Y(_07166_));
 sky130_fd_sc_hd__a21oi_1 _23817_ (.A1(_06985_),
    .A2(_06986_),
    .B1(_06987_),
    .Y(_07167_));
 sky130_fd_sc_hd__o21ai_2 _23818_ (.A1(_07166_),
    .A2(_07167_),
    .B1(_06989_),
    .Y(_07168_));
 sky130_vsdinv _23819_ (.A(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__nand2_1 _23820_ (.A(_07165_),
    .B(_07169_),
    .Y(_07170_));
 sky130_fd_sc_hd__nand3_2 _23821_ (.A(_07163_),
    .B(_07164_),
    .C(_07168_),
    .Y(_07171_));
 sky130_fd_sc_hd__nand2_1 _23822_ (.A(_07170_),
    .B(_07171_),
    .Y(_07172_));
 sky130_fd_sc_hd__o21ai_1 _23823_ (.A1(_06998_),
    .A2(_07006_),
    .B1(_06997_),
    .Y(_07173_));
 sky130_fd_sc_hd__xnor2_1 _23824_ (.A(_07172_),
    .B(_07173_),
    .Y(_02644_));
 sky130_fd_sc_hd__nand2_2 _23825_ (.A(_07157_),
    .B(_07149_),
    .Y(_07174_));
 sky130_fd_sc_hd__a31oi_4 _23826_ (.A1(_07063_),
    .A2(_07064_),
    .A3(_07139_),
    .B1(_07137_),
    .Y(_07175_));
 sky130_fd_sc_hd__a21o_1 _23827_ (.A1(_07010_),
    .A2(_07019_),
    .B1(_07021_),
    .X(_07176_));
 sky130_fd_sc_hd__or2b_1 _23828_ (.A(_07076_),
    .B_N(_07069_),
    .X(_07177_));
 sky130_fd_sc_hd__a21o_1 _23829_ (.A1(_06858_),
    .A2(_06860_),
    .B1(_07075_),
    .X(_07178_));
 sky130_fd_sc_hd__nand2_1 _23830_ (.A(_07177_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__nand3b_2 _23831_ (.A_N(_07014_),
    .B(_05127_),
    .C(_06285_),
    .Y(_07180_));
 sky130_fd_sc_hd__o31a_4 _23832_ (.A1(_14070_),
    .A2(_06293_),
    .A3(_07016_),
    .B1(_07180_),
    .X(_07181_));
 sky130_fd_sc_hd__nand3b_1 _23833_ (.A_N(_07066_),
    .B(_05879_),
    .C(_05610_),
    .Y(_07182_));
 sky130_fd_sc_hd__o31a_4 _23834_ (.A1(_05878_),
    .A2(_14365_),
    .A3(_07068_),
    .B1(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__and2_2 _23835_ (.A(_04996_),
    .B(_14337_),
    .X(_07184_));
 sky130_fd_sc_hd__nand2_2 _23836_ (.A(_05162_),
    .B(_14344_),
    .Y(_07185_));
 sky130_fd_sc_hd__and2_1 _23837_ (.A(_05129_),
    .B(\pcpi_mul.rs1[18] ),
    .X(_07186_));
 sky130_fd_sc_hd__xor2_4 _23838_ (.A(_07185_),
    .B(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__xor2_4 _23839_ (.A(_07184_),
    .B(_07187_),
    .X(_07188_));
 sky130_fd_sc_hd__xnor2_2 _23840_ (.A(_07183_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__xor2_2 _23841_ (.A(_07181_),
    .B(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__xnor2_1 _23842_ (.A(_07179_),
    .B(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__nor2_1 _23843_ (.A(_07012_),
    .B(_07017_),
    .Y(_07192_));
 sky130_fd_sc_hd__o21ba_1 _23844_ (.A1(_07011_),
    .A2(_07018_),
    .B1_N(_07192_),
    .X(_07193_));
 sky130_fd_sc_hd__nand2_1 _23845_ (.A(_07191_),
    .B(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__nor2_1 _23846_ (.A(_07193_),
    .B(_07191_),
    .Y(_07195_));
 sky130_vsdinv _23847_ (.A(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__and3_1 _23848_ (.A(_07176_),
    .B(_07194_),
    .C(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__clkbuf_4 _23849_ (.A(_06957_),
    .X(_07198_));
 sky130_fd_sc_hd__buf_6 _23850_ (.A(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__nor3_4 _23851_ (.A(_06433_),
    .B(_14329_),
    .C(_07041_),
    .Y(_07200_));
 sky130_fd_sc_hd__a41oi_4 _23852_ (.A1(_05298_),
    .A2(_04879_),
    .A3(_07199_),
    .A4(_07028_),
    .B1(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__a21oi_1 _23853_ (.A1(_06954_),
    .A2(_06958_),
    .B1(_07051_),
    .Y(_07202_));
 sky130_fd_sc_hd__o21bai_4 _23854_ (.A1(_07042_),
    .A2(_07052_),
    .B1_N(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__buf_2 _23855_ (.A(\pcpi_mul.rs1[23] ),
    .X(_07204_));
 sky130_fd_sc_hd__clkbuf_4 _23856_ (.A(_07204_),
    .X(_07205_));
 sky130_fd_sc_hd__buf_4 _23857_ (.A(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__and2_2 _23858_ (.A(_04932_),
    .B(_07206_),
    .X(_07207_));
 sky130_fd_sc_hd__nand2_2 _23859_ (.A(_04884_),
    .B(_07039_),
    .Y(_07208_));
 sky130_fd_sc_hd__buf_4 _23860_ (.A(\pcpi_mul.rs1[25] ),
    .X(_07209_));
 sky130_fd_sc_hd__buf_2 _23861_ (.A(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__nand2_2 _23862_ (.A(_04876_),
    .B(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__xnor2_4 _23863_ (.A(_07208_),
    .B(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__xor2_4 _23864_ (.A(_07207_),
    .B(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__buf_6 _23865_ (.A(_14332_),
    .X(_07214_));
 sky130_fd_sc_hd__a2bb2oi_4 _23866_ (.A1_N(_07214_),
    .A2_N(_07047_),
    .B1(_07045_),
    .B2(_07049_),
    .Y(_07215_));
 sky130_fd_sc_hd__clkbuf_4 _23867_ (.A(\pcpi_mul.rs1[26] ),
    .X(_07216_));
 sky130_fd_sc_hd__and2_2 _23868_ (.A(_04713_),
    .B(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__nand2_2 _23869_ (.A(_04924_),
    .B(_14325_),
    .Y(_07218_));
 sky130_fd_sc_hd__and2_1 _23870_ (.A(_14073_),
    .B(\pcpi_mul.rs1[21] ),
    .X(_07219_));
 sky130_fd_sc_hd__xor2_4 _23871_ (.A(_07218_),
    .B(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__xor2_4 _23872_ (.A(_07217_),
    .B(_07220_),
    .X(_07221_));
 sky130_fd_sc_hd__xnor2_4 _23873_ (.A(_07215_),
    .B(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__xor2_4 _23874_ (.A(_07213_),
    .B(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__xnor2_4 _23875_ (.A(_07203_),
    .B(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__xor2_4 _23876_ (.A(_07201_),
    .B(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__a21oi_2 _23877_ (.A1(_07194_),
    .A2(_07196_),
    .B1(_07176_),
    .Y(_07226_));
 sky130_vsdinv _23878_ (.A(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__nand3b_4 _23879_ (.A_N(_07197_),
    .B(_07225_),
    .C(_07227_),
    .Y(_07228_));
 sky130_fd_sc_hd__o21bai_2 _23880_ (.A1(_07226_),
    .A2(_07197_),
    .B1_N(_07225_),
    .Y(_07229_));
 sky130_fd_sc_hd__a21o_1 _23881_ (.A1(_07097_),
    .A2(_07098_),
    .B1(_07094_),
    .X(_07230_));
 sky130_fd_sc_hd__a21o_1 _23882_ (.A1(_07228_),
    .A2(_07229_),
    .B1(_07230_),
    .X(_07231_));
 sky130_fd_sc_hd__nand3_4 _23883_ (.A(_07228_),
    .B(_07230_),
    .C(_07229_),
    .Y(_07232_));
 sky130_fd_sc_hd__nor2_1 _23884_ (.A(_07026_),
    .B(_07056_),
    .Y(_07233_));
 sky130_vsdinv _23885_ (.A(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__a21oi_1 _23886_ (.A1(_07231_),
    .A2(_07232_),
    .B1(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__nand3_4 _23887_ (.A(_07231_),
    .B(_07234_),
    .C(_07232_),
    .Y(_07236_));
 sky130_fd_sc_hd__and2b_1 _23888_ (.A_N(_07235_),
    .B(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__a31oi_2 _23889_ (.A1(_07099_),
    .A2(_07133_),
    .A3(_07100_),
    .B1(_07131_),
    .Y(_07238_));
 sky130_fd_sc_hd__nor2_1 _23890_ (.A(_07122_),
    .B(_07124_),
    .Y(_07239_));
 sky130_fd_sc_hd__o21bai_1 _23891_ (.A1(_07117_),
    .A2(_07125_),
    .B1_N(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__and2_2 _23892_ (.A(_06060_),
    .B(_05875_),
    .X(_07241_));
 sky130_fd_sc_hd__nand2_2 _23893_ (.A(_14013_),
    .B(_05586_),
    .Y(_07242_));
 sky130_fd_sc_hd__and2_1 _23894_ (.A(_14008_),
    .B(_05089_),
    .X(_07243_));
 sky130_fd_sc_hd__xor2_4 _23895_ (.A(_07242_),
    .B(_07243_),
    .X(_07244_));
 sky130_fd_sc_hd__xor2_4 _23896_ (.A(_07241_),
    .B(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__buf_4 _23897_ (.A(_06744_),
    .X(_07246_));
 sky130_fd_sc_hd__buf_6 _23898_ (.A(_07246_),
    .X(_07247_));
 sky130_fd_sc_hd__nand3b_1 _23899_ (.A_N(_07119_),
    .B(_07247_),
    .C(_04937_),
    .Y(_07248_));
 sky130_fd_sc_hd__o31a_2 _23900_ (.A1(_07123_),
    .A2(_14434_),
    .A3(_07121_),
    .B1(_07248_),
    .X(_07249_));
 sky130_fd_sc_hd__and2_2 _23901_ (.A(_06470_),
    .B(_04978_),
    .X(_07250_));
 sky130_fd_sc_hd__nand2_2 _23902_ (.A(\pcpi_mul.rs2[22] ),
    .B(_04926_),
    .Y(_07251_));
 sky130_fd_sc_hd__and2_2 _23903_ (.A(\pcpi_mul.rs2[23] ),
    .B(\pcpi_mul.rs1[3] ),
    .X(_07252_));
 sky130_fd_sc_hd__xor2_4 _23904_ (.A(_07251_),
    .B(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__xor2_4 _23905_ (.A(_07250_),
    .B(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__xnor2_2 _23906_ (.A(_07249_),
    .B(_07254_),
    .Y(_07255_));
 sky130_fd_sc_hd__xor2_2 _23907_ (.A(_07245_),
    .B(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__xor2_1 _23908_ (.A(_07240_),
    .B(_07256_),
    .X(_07257_));
 sky130_fd_sc_hd__nor2_1 _23909_ (.A(_07105_),
    .B(_07108_),
    .Y(_07258_));
 sky130_vsdinv _23910_ (.A(_07258_),
    .Y(_07259_));
 sky130_fd_sc_hd__nand2_2 _23911_ (.A(_07106_),
    .B(_04937_),
    .Y(_07260_));
 sky130_fd_sc_hd__buf_2 _23912_ (.A(\pcpi_mul.rs2[26] ),
    .X(_07261_));
 sky130_fd_sc_hd__clkbuf_4 _23913_ (.A(_07261_),
    .X(_07262_));
 sky130_fd_sc_hd__nand3_4 _23914_ (.A(_07262_),
    .B(_07102_),
    .C(_04907_),
    .Y(_07263_));
 sky130_fd_sc_hd__clkbuf_4 _23915_ (.A(\pcpi_mul.rs2[26] ),
    .X(_07264_));
 sky130_fd_sc_hd__clkbuf_4 _23916_ (.A(_07101_),
    .X(_07265_));
 sky130_fd_sc_hd__a22o_1 _23917_ (.A1(_07264_),
    .A2(_05533_),
    .B1(_07265_),
    .B2(_14448_),
    .X(_07266_));
 sky130_fd_sc_hd__o21ai_2 _23918_ (.A1(_14452_),
    .A2(_07263_),
    .B1(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__xnor2_2 _23919_ (.A(_07260_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__xor2_1 _23920_ (.A(_07259_),
    .B(_07268_),
    .X(_07269_));
 sky130_fd_sc_hd__and2_1 _23921_ (.A(_07257_),
    .B(_07269_),
    .X(_07270_));
 sky130_vsdinv _23922_ (.A(_07128_),
    .Y(_07271_));
 sky130_fd_sc_hd__or2_2 _23923_ (.A(_07269_),
    .B(_07257_),
    .X(_07272_));
 sky130_fd_sc_hd__nor3b_4 _23924_ (.A(_07270_),
    .B(_07271_),
    .C_N(_07272_),
    .Y(_07273_));
 sky130_vsdinv _23925_ (.A(_07270_),
    .Y(_07274_));
 sky130_fd_sc_hd__a21oi_4 _23926_ (.A1(_07274_),
    .A2(_07272_),
    .B1(_07128_),
    .Y(_07275_));
 sky130_fd_sc_hd__and2_2 _23927_ (.A(_05720_),
    .B(_05913_),
    .X(_07276_));
 sky130_fd_sc_hd__nand2_2 _23928_ (.A(_14053_),
    .B(_05776_),
    .Y(_07277_));
 sky130_fd_sc_hd__and2_1 _23929_ (.A(_05357_),
    .B(_14370_),
    .X(_07278_));
 sky130_fd_sc_hd__xor2_4 _23930_ (.A(_07277_),
    .B(_07278_),
    .X(_07279_));
 sky130_fd_sc_hd__xnor2_4 _23931_ (.A(_07276_),
    .B(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__buf_4 _23932_ (.A(_05635_),
    .X(_07281_));
 sky130_fd_sc_hd__nand3b_1 _23933_ (.A_N(_07072_),
    .B(_07281_),
    .C(_05413_),
    .Y(_07282_));
 sky130_fd_sc_hd__o31a_2 _23934_ (.A1(_06207_),
    .A2(_14383_),
    .A3(_07074_),
    .B1(_07282_),
    .X(_07283_));
 sky130_fd_sc_hd__and2_2 _23935_ (.A(_05440_),
    .B(_06412_),
    .X(_07284_));
 sky130_fd_sc_hd__nand2_2 _23936_ (.A(_06855_),
    .B(_14381_),
    .Y(_07285_));
 sky130_fd_sc_hd__and2_1 _23937_ (.A(_05634_),
    .B(\pcpi_mul.rs1[12] ),
    .X(_07286_));
 sky130_fd_sc_hd__xor2_4 _23938_ (.A(_07285_),
    .B(_07286_),
    .X(_07287_));
 sky130_fd_sc_hd__xor2_4 _23939_ (.A(_07284_),
    .B(_07287_),
    .X(_07288_));
 sky130_fd_sc_hd__xnor2_1 _23940_ (.A(_07283_),
    .B(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__xnor2_1 _23941_ (.A(_07280_),
    .B(_07289_),
    .Y(_07290_));
 sky130_vsdinv _23942_ (.A(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__nor2_1 _23943_ (.A(_07082_),
    .B(_07087_),
    .Y(_07292_));
 sky130_fd_sc_hd__o21bai_1 _23944_ (.A1(_07081_),
    .A2(_07088_),
    .B1_N(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__buf_4 _23945_ (.A(_14023_),
    .X(_07294_));
 sky130_fd_sc_hd__buf_6 _23946_ (.A(_07294_),
    .X(_07295_));
 sky130_fd_sc_hd__nand3b_1 _23947_ (.A_N(_07084_),
    .B(_07295_),
    .C(_05229_),
    .Y(_07296_));
 sky130_fd_sc_hd__o31a_2 _23948_ (.A1(_14033_),
    .A2(_14401_),
    .A3(_07086_),
    .B1(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__nand3b_1 _23949_ (.A_N(_07114_),
    .B(_06895_),
    .C(_05039_),
    .Y(_07298_));
 sky130_fd_sc_hd__o31a_2 _23950_ (.A1(_14018_),
    .A2(_05115_),
    .A3(_07116_),
    .B1(_07298_),
    .X(_07299_));
 sky130_fd_sc_hd__and2_2 _23951_ (.A(_05716_),
    .B(_05321_),
    .X(_07300_));
 sky130_fd_sc_hd__nand2_2 _23952_ (.A(_06351_),
    .B(_05613_),
    .Y(_07301_));
 sky130_fd_sc_hd__and2_1 _23953_ (.A(_06485_),
    .B(_05180_),
    .X(_07302_));
 sky130_fd_sc_hd__xor2_4 _23954_ (.A(_07301_),
    .B(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__xor2_4 _23955_ (.A(_07300_),
    .B(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__xnor2_2 _23956_ (.A(_07299_),
    .B(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__xor2_2 _23957_ (.A(_07297_),
    .B(_07305_),
    .X(_07306_));
 sky130_fd_sc_hd__xnor2_1 _23958_ (.A(_07293_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__nor2_1 _23959_ (.A(_07291_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__and2_1 _23960_ (.A(_07126_),
    .B(_07112_),
    .X(_07309_));
 sky130_fd_sc_hd__nand2_1 _23961_ (.A(_07307_),
    .B(_07291_),
    .Y(_07310_));
 sky130_fd_sc_hd__and3b_1 _23962_ (.A_N(_07308_),
    .B(_07309_),
    .C(_07310_),
    .X(_07311_));
 sky130_vsdinv _23963_ (.A(_07311_),
    .Y(_07312_));
 sky130_vsdinv _23964_ (.A(_07308_),
    .Y(_07313_));
 sky130_fd_sc_hd__a21o_2 _23965_ (.A1(_07313_),
    .A2(_07310_),
    .B1(_07309_),
    .X(_07314_));
 sky130_fd_sc_hd__a21o_2 _23966_ (.A1(_07089_),
    .A2(_07080_),
    .B1(_07091_),
    .X(_07315_));
 sky130_fd_sc_hd__a21oi_4 _23967_ (.A1(_07312_),
    .A2(_07314_),
    .B1(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__nand3b_4 _23968_ (.A_N(_07311_),
    .B(_07315_),
    .C(_07314_),
    .Y(_07317_));
 sky130_vsdinv _23969_ (.A(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__o22ai_4 _23970_ (.A1(_07273_),
    .A2(_07275_),
    .B1(_07316_),
    .B2(_07318_),
    .Y(_07319_));
 sky130_fd_sc_hd__nor2_2 _23971_ (.A(_07273_),
    .B(_07275_),
    .Y(_07320_));
 sky130_fd_sc_hd__nand3b_4 _23972_ (.A_N(_07316_),
    .B(_07317_),
    .C(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__nand3b_4 _23973_ (.A_N(_07238_),
    .B(_07319_),
    .C(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__a21bo_2 _23974_ (.A1(_07321_),
    .A2(_07319_),
    .B1_N(_07238_),
    .X(_07323_));
 sky130_fd_sc_hd__nand3_4 _23975_ (.A(_07237_),
    .B(_07322_),
    .C(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__a21boi_4 _23976_ (.A1(_07319_),
    .A2(_07321_),
    .B1_N(_07238_),
    .Y(_07325_));
 sky130_vsdinv _23977_ (.A(_07322_),
    .Y(_07326_));
 sky130_vsdinv _23978_ (.A(_07235_),
    .Y(_07327_));
 sky130_fd_sc_hd__nand2_1 _23979_ (.A(_07327_),
    .B(_07236_),
    .Y(_07328_));
 sky130_fd_sc_hd__o21ai_2 _23980_ (.A1(_07325_),
    .A2(_07326_),
    .B1(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__nand3b_4 _23981_ (.A_N(_07175_),
    .B(_07324_),
    .C(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand2_1 _23982_ (.A(_07324_),
    .B(_07329_),
    .Y(_07331_));
 sky130_fd_sc_hd__nand2_2 _23983_ (.A(_07331_),
    .B(_07175_),
    .Y(_07332_));
 sky130_fd_sc_hd__nor2_2 _23984_ (.A(_07030_),
    .B(_07054_),
    .Y(_07333_));
 sky130_fd_sc_hd__a21oi_4 _23985_ (.A1(_07053_),
    .A2(_07032_),
    .B1(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__a21oi_4 _23986_ (.A1(_07064_),
    .A2(_07061_),
    .B1(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__and3_1 _23987_ (.A(_07064_),
    .B(_07061_),
    .C(_07334_),
    .X(_07336_));
 sky130_fd_sc_hd__o2bb2ai_2 _23988_ (.A1_N(_07330_),
    .A2_N(_07332_),
    .B1(_07335_),
    .B2(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__nor2_2 _23989_ (.A(_07335_),
    .B(_07336_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand3_4 _23990_ (.A(_07332_),
    .B(_07330_),
    .C(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__nand3_4 _23991_ (.A(_07174_),
    .B(_07337_),
    .C(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand2_1 _23992_ (.A(_07337_),
    .B(_07339_),
    .Y(_07341_));
 sky130_fd_sc_hd__a21boi_1 _23993_ (.A1(_07146_),
    .A2(_07154_),
    .B1_N(_07149_),
    .Y(_07342_));
 sky130_fd_sc_hd__nand2_1 _23994_ (.A(_07341_),
    .B(_07342_),
    .Y(_07343_));
 sky130_fd_sc_hd__o2bb2ai_1 _23995_ (.A1_N(_07340_),
    .A2_N(_07343_),
    .B1(_07153_),
    .B2(_07152_),
    .Y(_07344_));
 sky130_fd_sc_hd__nor2_2 _23996_ (.A(_07152_),
    .B(_07153_),
    .Y(_07345_));
 sky130_fd_sc_hd__nand3_2 _23997_ (.A(_07343_),
    .B(_07345_),
    .C(_07340_),
    .Y(_07346_));
 sky130_vsdinv _23998_ (.A(_07162_),
    .Y(_07347_));
 sky130_fd_sc_hd__o21ai_1 _23999_ (.A1(_07347_),
    .A2(_07159_),
    .B1(_07160_),
    .Y(_07348_));
 sky130_fd_sc_hd__a21oi_1 _24000_ (.A1(_07344_),
    .A2(_07346_),
    .B1(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand3_1 _24001_ (.A(_07344_),
    .B(_07346_),
    .C(_07348_),
    .Y(_07350_));
 sky130_vsdinv _24002_ (.A(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__nor2_2 _24003_ (.A(_07349_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__and2_1 _24004_ (.A(_05868_),
    .B(_07000_),
    .X(_07353_));
 sky130_fd_sc_hd__o21bai_1 _24005_ (.A1(_07005_),
    .A2(_07353_),
    .B1_N(_07172_),
    .Y(_07354_));
 sky130_fd_sc_hd__a21oi_1 _24006_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07168_),
    .Y(_07355_));
 sky130_fd_sc_hd__a21oi_2 _24007_ (.A1(_06997_),
    .A2(_07171_),
    .B1(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__o21bai_1 _24008_ (.A1(_06998_),
    .A2(_07354_),
    .B1_N(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__xor2_1 _24009_ (.A(_07352_),
    .B(_07357_),
    .X(_02645_));
 sky130_fd_sc_hd__buf_2 _24010_ (.A(\pcpi_mul.rs2[27] ),
    .X(_07358_));
 sky130_fd_sc_hd__buf_6 _24011_ (.A(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__buf_6 _24012_ (.A(_07359_),
    .X(_07360_));
 sky130_fd_sc_hd__nand2_8 _24013_ (.A(_07360_),
    .B(_04719_),
    .Y(_07361_));
 sky130_fd_sc_hd__o22a_4 _24014_ (.A1(_14453_),
    .A2(_07263_),
    .B1(_07260_),
    .B2(_07267_),
    .X(_07362_));
 sky130_fd_sc_hd__and2_2 _24015_ (.A(_06887_),
    .B(_04898_),
    .X(_07363_));
 sky130_fd_sc_hd__nand2_2 _24016_ (.A(_07261_),
    .B(_04906_),
    .Y(_07364_));
 sky130_fd_sc_hd__nand2_2 _24017_ (.A(_07101_),
    .B(_04889_),
    .Y(_07365_));
 sky130_fd_sc_hd__xnor2_4 _24018_ (.A(_07364_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__xor2_4 _24019_ (.A(_07363_),
    .B(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__xnor2_4 _24020_ (.A(_07362_),
    .B(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__xor2_4 _24021_ (.A(_07361_),
    .B(_07368_),
    .X(_07369_));
 sky130_fd_sc_hd__nor2_1 _24022_ (.A(_07249_),
    .B(_07254_),
    .Y(_07370_));
 sky130_fd_sc_hd__o21ba_2 _24023_ (.A1(_07245_),
    .A2(_07255_),
    .B1_N(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__or2b_4 _24024_ (.A(_07268_),
    .B_N(_07258_),
    .X(_07372_));
 sky130_fd_sc_hd__and2_1 _24025_ (.A(_06319_),
    .B(_05308_),
    .X(_07373_));
 sky130_fd_sc_hd__nand3_4 _24026_ (.A(_06321_),
    .B(_06737_),
    .C(_05429_),
    .Y(_07374_));
 sky130_fd_sc_hd__a22o_1 _24027_ (.A1(_06321_),
    .A2(_05047_),
    .B1(_06737_),
    .B2(_05105_),
    .X(_07375_));
 sky130_fd_sc_hd__o21ai_1 _24028_ (.A1(_05998_),
    .A2(_07374_),
    .B1(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__xnor2_1 _24029_ (.A(_07373_),
    .B(_07376_),
    .Y(_07377_));
 sky130_vsdinv _24030_ (.A(_07377_),
    .Y(_07378_));
 sky130_fd_sc_hd__nand3b_1 _24031_ (.A_N(_07251_),
    .B(_07246_),
    .C(_04898_),
    .Y(_07379_));
 sky130_fd_sc_hd__o31a_2 _24032_ (.A1(_14005_),
    .A2(_14428_),
    .A3(_07253_),
    .B1(_07379_),
    .X(_07380_));
 sky130_fd_sc_hd__and2_2 _24033_ (.A(_06469_),
    .B(_05098_),
    .X(_07381_));
 sky130_fd_sc_hd__nand2_2 _24034_ (.A(\pcpi_mul.rs2[22] ),
    .B(_14426_),
    .Y(_07382_));
 sky130_fd_sc_hd__and2_2 _24035_ (.A(\pcpi_mul.rs2[23] ),
    .B(\pcpi_mul.rs1[4] ),
    .X(_07383_));
 sky130_fd_sc_hd__xor2_4 _24036_ (.A(_07382_),
    .B(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__xor2_4 _24037_ (.A(_07381_),
    .B(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__xnor2_4 _24038_ (.A(_07380_),
    .B(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__xor2_4 _24039_ (.A(_07378_),
    .B(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__xor2_4 _24040_ (.A(_07372_),
    .B(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__xor2_4 _24041_ (.A(_07371_),
    .B(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__nor2_2 _24042_ (.A(_07369_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__and2_2 _24043_ (.A(_07389_),
    .B(_07369_),
    .X(_07391_));
 sky130_fd_sc_hd__nor3_4 _24044_ (.A(_07274_),
    .B(_07390_),
    .C(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__o21a_1 _24045_ (.A1(_07390_),
    .A2(_07391_),
    .B1(_07274_),
    .X(_07393_));
 sky130_fd_sc_hd__and2_2 _24046_ (.A(_05205_),
    .B(_06288_),
    .X(_07394_));
 sky130_fd_sc_hd__nand2_2 _24047_ (.A(_14053_),
    .B(_14357_),
    .Y(_07395_));
 sky130_fd_sc_hd__and2_1 _24048_ (.A(\pcpi_mul.rs2[11] ),
    .B(\pcpi_mul.rs1[16] ),
    .X(_07396_));
 sky130_fd_sc_hd__xor2_4 _24049_ (.A(_07395_),
    .B(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__xnor2_4 _24050_ (.A(_07394_),
    .B(_07397_),
    .Y(_07398_));
 sky130_fd_sc_hd__nand3b_2 _24051_ (.A_N(_07285_),
    .B(_14037_),
    .C(_05423_),
    .Y(_07399_));
 sky130_fd_sc_hd__o31a_4 _24052_ (.A1(_14046_),
    .A2(_06264_),
    .A3(_07287_),
    .B1(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__and2_2 _24053_ (.A(_05727_),
    .B(_05698_),
    .X(_07401_));
 sky130_fd_sc_hd__nand2_2 _24054_ (.A(_06855_),
    .B(\pcpi_mul.rs1[14] ),
    .Y(_07402_));
 sky130_fd_sc_hd__and2_1 _24055_ (.A(_14035_),
    .B(_14381_),
    .X(_07403_));
 sky130_fd_sc_hd__xor2_4 _24056_ (.A(_07402_),
    .B(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__xor2_4 _24057_ (.A(_07401_),
    .B(_07404_),
    .X(_07405_));
 sky130_fd_sc_hd__xnor2_4 _24058_ (.A(_07400_),
    .B(_07405_),
    .Y(_07406_));
 sky130_fd_sc_hd__xnor2_4 _24059_ (.A(_07398_),
    .B(_07406_),
    .Y(_07407_));
 sky130_vsdinv _24060_ (.A(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__nor2_1 _24061_ (.A(_07299_),
    .B(_07304_),
    .Y(_07409_));
 sky130_fd_sc_hd__o21bai_1 _24062_ (.A1(_07297_),
    .A2(_07305_),
    .B1_N(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__nand3b_1 _24063_ (.A_N(_07301_),
    .B(_07295_),
    .C(_05301_),
    .Y(_07411_));
 sky130_fd_sc_hd__o31a_2 _24064_ (.A1(_14033_),
    .A2(_14395_),
    .A3(_07303_),
    .B1(_07411_),
    .X(_07412_));
 sky130_fd_sc_hd__nand3b_1 _24065_ (.A_N(_07242_),
    .B(_06322_),
    .C(_05099_),
    .Y(_07413_));
 sky130_fd_sc_hd__o31a_1 _24066_ (.A1(_14018_),
    .A2(_14411_),
    .A3(_07244_),
    .B1(_07413_),
    .X(_07414_));
 sky130_fd_sc_hd__and2_2 _24067_ (.A(\pcpi_mul.rs2[15] ),
    .B(_06002_),
    .X(_07415_));
 sky130_fd_sc_hd__nand2_2 _24068_ (.A(_06070_),
    .B(_05320_),
    .Y(_07416_));
 sky130_fd_sc_hd__and2_1 _24069_ (.A(_14022_),
    .B(_14398_),
    .X(_07417_));
 sky130_fd_sc_hd__xor2_4 _24070_ (.A(_07416_),
    .B(_07417_),
    .X(_07418_));
 sky130_fd_sc_hd__xor2_4 _24071_ (.A(_07415_),
    .B(_07418_),
    .X(_07419_));
 sky130_fd_sc_hd__xnor2_2 _24072_ (.A(_07414_),
    .B(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__xor2_2 _24073_ (.A(_07412_),
    .B(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__xnor2_1 _24074_ (.A(_07410_),
    .B(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__nor2_1 _24075_ (.A(_07408_),
    .B(_07422_),
    .Y(_07423_));
 sky130_vsdinv _24076_ (.A(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__nand2_1 _24077_ (.A(_07422_),
    .B(_07408_),
    .Y(_07425_));
 sky130_fd_sc_hd__and2_1 _24078_ (.A(_07256_),
    .B(_07240_),
    .X(_07426_));
 sky130_fd_sc_hd__a21oi_2 _24079_ (.A1(_07424_),
    .A2(_07425_),
    .B1(_07426_),
    .Y(_07427_));
 sky130_fd_sc_hd__and3b_1 _24080_ (.A_N(_07423_),
    .B(_07426_),
    .C(_07425_),
    .X(_07428_));
 sky130_vsdinv _24081_ (.A(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__nand2_1 _24082_ (.A(_07306_),
    .B(_07293_),
    .Y(_07430_));
 sky130_fd_sc_hd__o21a_1 _24083_ (.A1(_07291_),
    .A2(_07307_),
    .B1(_07430_),
    .X(_07431_));
 sky130_vsdinv _24084_ (.A(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__nand3b_1 _24085_ (.A_N(_07427_),
    .B(_07429_),
    .C(_07432_),
    .Y(_07433_));
 sky130_fd_sc_hd__o21bai_1 _24086_ (.A1(_07427_),
    .A2(_07428_),
    .B1_N(_07432_),
    .Y(_07434_));
 sky130_fd_sc_hd__nand2_2 _24087_ (.A(_07433_),
    .B(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__o21a_2 _24088_ (.A1(_07392_),
    .A2(_07393_),
    .B1(_07435_),
    .X(_07436_));
 sky130_fd_sc_hd__nor3_4 _24089_ (.A(_07392_),
    .B(_07393_),
    .C(_07435_),
    .Y(_07437_));
 sky130_vsdinv _24090_ (.A(_07273_),
    .Y(_07438_));
 sky130_fd_sc_hd__o211ai_4 _24091_ (.A1(_07436_),
    .A2(_07437_),
    .B1(_07438_),
    .C1(_07321_),
    .Y(_07439_));
 sky130_vsdinv _24092_ (.A(_07436_),
    .Y(_07440_));
 sky130_fd_sc_hd__nand2_1 _24093_ (.A(_07321_),
    .B(_07438_),
    .Y(_07441_));
 sky130_fd_sc_hd__nand3b_4 _24094_ (.A_N(_07437_),
    .B(_07440_),
    .C(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__and2_1 _24095_ (.A(_07190_),
    .B(_07179_),
    .X(_07443_));
 sky130_fd_sc_hd__nand3b_1 _24096_ (.A_N(_07185_),
    .B(_05577_),
    .C(_06280_),
    .Y(_07444_));
 sky130_fd_sc_hd__o31a_2 _24097_ (.A1(_05576_),
    .A2(_14341_),
    .A3(_07187_),
    .B1(_07444_),
    .X(_07445_));
 sky130_fd_sc_hd__nand3b_1 _24098_ (.A_N(_07277_),
    .B(_05359_),
    .C(_05769_),
    .Y(_07446_));
 sky130_fd_sc_hd__o31a_2 _24099_ (.A1(_05878_),
    .A2(_14359_),
    .A3(_07279_),
    .B1(_07446_),
    .X(_07447_));
 sky130_fd_sc_hd__and2_2 _24100_ (.A(_05483_),
    .B(_14331_),
    .X(_07448_));
 sky130_fd_sc_hd__nand2_2 _24101_ (.A(_05063_),
    .B(_14337_),
    .Y(_07449_));
 sky130_fd_sc_hd__and2_1 _24102_ (.A(_05130_),
    .B(_14344_),
    .X(_07450_));
 sky130_fd_sc_hd__xor2_4 _24103_ (.A(_07449_),
    .B(_07450_),
    .X(_07451_));
 sky130_fd_sc_hd__xor2_4 _24104_ (.A(_07448_),
    .B(_07451_),
    .X(_07452_));
 sky130_fd_sc_hd__xnor2_4 _24105_ (.A(_07447_),
    .B(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__xor2_4 _24106_ (.A(_07445_),
    .B(_07453_),
    .X(_07454_));
 sky130_fd_sc_hd__or2b_1 _24107_ (.A(_07289_),
    .B_N(_07280_),
    .X(_07455_));
 sky130_fd_sc_hd__o21ai_2 _24108_ (.A1(_07288_),
    .A2(_07283_),
    .B1(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__xnor2_1 _24109_ (.A(_07454_),
    .B(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__nor2_1 _24110_ (.A(_07183_),
    .B(_07188_),
    .Y(_07458_));
 sky130_fd_sc_hd__o21ba_1 _24111_ (.A1(_07181_),
    .A2(_07189_),
    .B1_N(_07458_),
    .X(_07459_));
 sky130_fd_sc_hd__nand2_1 _24112_ (.A(_07457_),
    .B(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__nor2_1 _24113_ (.A(_07459_),
    .B(_07457_),
    .Y(_07461_));
 sky130_vsdinv _24114_ (.A(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__o211a_1 _24115_ (.A1(_07443_),
    .A2(_07195_),
    .B1(_07460_),
    .C1(_07462_),
    .X(_07463_));
 sky130_vsdinv _24116_ (.A(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__o21bai_1 _24117_ (.A1(_07193_),
    .A2(_07191_),
    .B1_N(_07443_),
    .Y(_07465_));
 sky130_fd_sc_hd__a21o_1 _24118_ (.A1(_07462_),
    .A2(_07460_),
    .B1(_07465_),
    .X(_07466_));
 sky130_fd_sc_hd__clkbuf_4 _24119_ (.A(_07044_),
    .X(_07467_));
 sky130_fd_sc_hd__buf_6 _24120_ (.A(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__nor3_4 _24121_ (.A(_14087_),
    .B(_14322_),
    .C(_07212_),
    .Y(_07469_));
 sky130_fd_sc_hd__a41oi_4 _24122_ (.A1(_05403_),
    .A2(_05300_),
    .A3(_07468_),
    .A4(_07199_),
    .B1(_07469_),
    .Y(_07470_));
 sky130_fd_sc_hd__nor2_1 _24123_ (.A(_07215_),
    .B(_07221_),
    .Y(_07471_));
 sky130_fd_sc_hd__o21bai_4 _24124_ (.A1(_07213_),
    .A2(_07222_),
    .B1_N(_07471_),
    .Y(_07472_));
 sky130_fd_sc_hd__buf_2 _24125_ (.A(_07039_),
    .X(_07473_));
 sky130_fd_sc_hd__and2_2 _24126_ (.A(_14083_),
    .B(_07473_),
    .X(_07474_));
 sky130_fd_sc_hd__nand2_2 _24127_ (.A(_04905_),
    .B(_07210_),
    .Y(_07475_));
 sky130_fd_sc_hd__buf_2 _24128_ (.A(\pcpi_mul.rs1[26] ),
    .X(_07476_));
 sky130_fd_sc_hd__clkbuf_4 _24129_ (.A(_07476_),
    .X(_07477_));
 sky130_fd_sc_hd__nand2_2 _24130_ (.A(_04910_),
    .B(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__xnor2_4 _24131_ (.A(_07475_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__xor2_4 _24132_ (.A(_07474_),
    .B(_07479_),
    .X(_07480_));
 sky130_fd_sc_hd__clkbuf_4 _24133_ (.A(_06450_),
    .X(_07481_));
 sky130_fd_sc_hd__nand3b_1 _24134_ (.A_N(_07218_),
    .B(_05420_),
    .C(_07481_),
    .Y(_07482_));
 sky130_fd_sc_hd__o31a_2 _24135_ (.A1(_05315_),
    .A2(_14304_),
    .A3(_07220_),
    .B1(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__clkbuf_2 _24136_ (.A(\pcpi_mul.rs1[27] ),
    .X(_07484_));
 sky130_fd_sc_hd__buf_2 _24137_ (.A(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__and2_2 _24138_ (.A(_05319_),
    .B(_07485_),
    .X(_07486_));
 sky130_fd_sc_hd__nand2_2 _24139_ (.A(_05324_),
    .B(_06777_),
    .Y(_07487_));
 sky130_fd_sc_hd__and2_1 _24140_ (.A(_05326_),
    .B(_06939_),
    .X(_07488_));
 sky130_fd_sc_hd__xor2_4 _24141_ (.A(_07487_),
    .B(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__xor2_4 _24142_ (.A(_07486_),
    .B(_07489_),
    .X(_07490_));
 sky130_fd_sc_hd__xnor2_4 _24143_ (.A(_07483_),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__xor2_4 _24144_ (.A(_07480_),
    .B(_07491_),
    .X(_07492_));
 sky130_fd_sc_hd__xnor2_4 _24145_ (.A(_07472_),
    .B(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__xor2_4 _24146_ (.A(_07470_),
    .B(_07493_),
    .X(_07494_));
 sky130_fd_sc_hd__a21o_1 _24147_ (.A1(_07464_),
    .A2(_07466_),
    .B1(_07494_),
    .X(_07495_));
 sky130_fd_sc_hd__nand3b_4 _24148_ (.A_N(_07463_),
    .B(_07494_),
    .C(_07466_),
    .Y(_07496_));
 sky130_fd_sc_hd__a21o_1 _24149_ (.A1(_07314_),
    .A2(_07315_),
    .B1(_07311_),
    .X(_07497_));
 sky130_fd_sc_hd__a21o_1 _24150_ (.A1(_07495_),
    .A2(_07496_),
    .B1(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__a21oi_1 _24151_ (.A1(_07227_),
    .A2(_07225_),
    .B1(_07197_),
    .Y(_07499_));
 sky130_vsdinv _24152_ (.A(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__nand3_4 _24153_ (.A(_07495_),
    .B(_07497_),
    .C(_07496_),
    .Y(_07501_));
 sky130_fd_sc_hd__nand3_1 _24154_ (.A(_07498_),
    .B(_07500_),
    .C(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__clkbuf_4 _24155_ (.A(_07502_),
    .X(_07503_));
 sky130_fd_sc_hd__a21o_2 _24156_ (.A1(_07498_),
    .A2(_07501_),
    .B1(_07500_),
    .X(_07504_));
 sky130_fd_sc_hd__a22oi_4 _24157_ (.A1(_07439_),
    .A2(_07442_),
    .B1(_07503_),
    .B2(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__nand2_1 _24158_ (.A(_07439_),
    .B(_07442_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand2_1 _24159_ (.A(_07504_),
    .B(_07503_),
    .Y(_07507_));
 sky130_fd_sc_hd__nor2_2 _24160_ (.A(_07506_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__a31oi_4 _24161_ (.A1(_07323_),
    .A2(_07327_),
    .A3(_07236_),
    .B1(_07326_),
    .Y(_07509_));
 sky130_fd_sc_hd__o21ai_4 _24162_ (.A1(_07505_),
    .A2(_07508_),
    .B1(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__o21bai_2 _24163_ (.A1(_07325_),
    .A2(_07328_),
    .B1_N(_07326_),
    .Y(_07511_));
 sky130_fd_sc_hd__a21oi_2 _24164_ (.A1(_07498_),
    .A2(_07501_),
    .B1(_07500_),
    .Y(_07512_));
 sky130_vsdinv _24165_ (.A(_07502_),
    .Y(_07513_));
 sky130_fd_sc_hd__nor2_1 _24166_ (.A(_07512_),
    .B(_07513_),
    .Y(_07514_));
 sky130_fd_sc_hd__nand3_2 _24167_ (.A(_07514_),
    .B(_07442_),
    .C(_07439_),
    .Y(_07515_));
 sky130_fd_sc_hd__o2bb2ai_2 _24168_ (.A1_N(_07442_),
    .A2_N(_07439_),
    .B1(_07512_),
    .B2(_07513_),
    .Y(_07516_));
 sky130_fd_sc_hd__nand3_4 _24169_ (.A(_07511_),
    .B(_07515_),
    .C(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__nand2_1 _24170_ (.A(_07510_),
    .B(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__nor2_1 _24171_ (.A(_07201_),
    .B(_07224_),
    .Y(_07519_));
 sky130_fd_sc_hd__a21o_4 _24172_ (.A1(_07223_),
    .A2(_07203_),
    .B1(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__nand2_2 _24173_ (.A(_07236_),
    .B(_07232_),
    .Y(_07521_));
 sky130_fd_sc_hd__xor2_4 _24174_ (.A(_07520_),
    .B(_07521_),
    .X(_07522_));
 sky130_vsdinv _24175_ (.A(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__nand2_2 _24176_ (.A(_07518_),
    .B(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__nand3_4 _24177_ (.A(_07510_),
    .B(_07522_),
    .C(_07517_),
    .Y(_07525_));
 sky130_fd_sc_hd__nand2_4 _24178_ (.A(_07339_),
    .B(_07330_),
    .Y(_07526_));
 sky130_fd_sc_hd__a21o_1 _24179_ (.A1(_07524_),
    .A2(_07525_),
    .B1(_07526_),
    .X(_07527_));
 sky130_fd_sc_hd__nand3_4 _24180_ (.A(_07526_),
    .B(_07524_),
    .C(_07525_),
    .Y(_07528_));
 sky130_fd_sc_hd__a21oi_1 _24181_ (.A1(_07527_),
    .A2(_07528_),
    .B1(_07335_),
    .Y(_07529_));
 sky130_vsdinv _24182_ (.A(_07335_),
    .Y(_07530_));
 sky130_fd_sc_hd__a21oi_4 _24183_ (.A1(_07524_),
    .A2(_07525_),
    .B1(_07526_),
    .Y(_07531_));
 sky130_fd_sc_hd__nor3b_2 _24184_ (.A(_07530_),
    .B(_07531_),
    .C_N(_07528_),
    .Y(_07532_));
 sky130_vsdinv _24185_ (.A(_07345_),
    .Y(_07533_));
 sky130_fd_sc_hd__a21oi_1 _24186_ (.A1(_07337_),
    .A2(_07339_),
    .B1(_07174_),
    .Y(_07534_));
 sky130_fd_sc_hd__o21ai_1 _24187_ (.A1(_07533_),
    .A2(_07534_),
    .B1(_07340_),
    .Y(_07535_));
 sky130_fd_sc_hd__o21bai_1 _24188_ (.A1(_07529_),
    .A2(_07532_),
    .B1_N(_07535_),
    .Y(_07536_));
 sky130_vsdinv _24189_ (.A(_07528_),
    .Y(_07537_));
 sky130_fd_sc_hd__o21bai_1 _24190_ (.A1(_07531_),
    .A2(_07537_),
    .B1_N(_07335_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand3_1 _24191_ (.A(_07527_),
    .B(_07335_),
    .C(_07528_),
    .Y(_07539_));
 sky130_fd_sc_hd__nand3_1 _24192_ (.A(_07538_),
    .B(_07539_),
    .C(_07535_),
    .Y(_07540_));
 sky130_fd_sc_hd__nand2_1 _24193_ (.A(_07536_),
    .B(_07540_),
    .Y(_07541_));
 sky130_fd_sc_hd__a21oi_1 _24194_ (.A1(_07343_),
    .A2(_07340_),
    .B1(_07345_),
    .Y(_07542_));
 sky130_vsdinv _24195_ (.A(_07346_),
    .Y(_07543_));
 sky130_fd_sc_hd__o21bai_1 _24196_ (.A1(_07542_),
    .A2(_07543_),
    .B1_N(_07348_),
    .Y(_07544_));
 sky130_fd_sc_hd__a21oi_1 _24197_ (.A1(_07357_),
    .A2(_07544_),
    .B1(_07351_),
    .Y(_07545_));
 sky130_fd_sc_hd__xor2_1 _24198_ (.A(_07541_),
    .B(_07545_),
    .X(_02646_));
 sky130_fd_sc_hd__nand3b_1 _24199_ (.A_N(_07449_),
    .B(_05577_),
    .C(_06584_),
    .Y(_07546_));
 sky130_fd_sc_hd__o31a_2 _24200_ (.A1(_05576_),
    .A2(_07214_),
    .A3(_07451_),
    .B1(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__nand3b_1 _24201_ (.A_N(_07395_),
    .B(_05361_),
    .C(_05777_),
    .Y(_07548_));
 sky130_fd_sc_hd__o31a_2 _24202_ (.A1(_05878_),
    .A2(_14352_),
    .A3(_07397_),
    .B1(_07548_),
    .X(_07549_));
 sky130_fd_sc_hd__and2_2 _24203_ (.A(_06001_),
    .B(_14325_),
    .X(_07550_));
 sky130_fd_sc_hd__nand2_2 _24204_ (.A(_05063_),
    .B(\pcpi_mul.rs1[21] ),
    .Y(_07551_));
 sky130_fd_sc_hd__and2_1 _24205_ (.A(_14061_),
    .B(_14337_),
    .X(_07552_));
 sky130_fd_sc_hd__xor2_4 _24206_ (.A(_07551_),
    .B(_07552_),
    .X(_07553_));
 sky130_fd_sc_hd__xor2_4 _24207_ (.A(_07550_),
    .B(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__xnor2_4 _24208_ (.A(_07549_),
    .B(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__xor2_4 _24209_ (.A(_07547_),
    .B(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__or2b_1 _24210_ (.A(_07406_),
    .B_N(_07398_),
    .X(_07557_));
 sky130_fd_sc_hd__o21ai_4 _24211_ (.A1(_07405_),
    .A2(_07400_),
    .B1(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__xnor2_1 _24212_ (.A(_07556_),
    .B(_07558_),
    .Y(_07559_));
 sky130_fd_sc_hd__nor2_1 _24213_ (.A(_07447_),
    .B(_07452_),
    .Y(_07560_));
 sky130_fd_sc_hd__o21ba_2 _24214_ (.A1(_07445_),
    .A2(_07453_),
    .B1_N(_07560_),
    .X(_07561_));
 sky130_fd_sc_hd__nand2_2 _24215_ (.A(_07559_),
    .B(_07561_),
    .Y(_07562_));
 sky130_fd_sc_hd__nor2_1 _24216_ (.A(_07561_),
    .B(_07559_),
    .Y(_07563_));
 sky130_vsdinv _24217_ (.A(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__a21o_1 _24218_ (.A1(_07456_),
    .A2(_07454_),
    .B1(_07461_),
    .X(_07565_));
 sky130_fd_sc_hd__a21o_1 _24219_ (.A1(_07562_),
    .A2(_07564_),
    .B1(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__nand3_4 _24220_ (.A(_07565_),
    .B(_07564_),
    .C(_07562_),
    .Y(_07567_));
 sky130_fd_sc_hd__buf_4 _24221_ (.A(\pcpi_mul.rs1[26] ),
    .X(_07568_));
 sky130_fd_sc_hd__clkbuf_4 _24222_ (.A(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__buf_4 _24223_ (.A(_07569_),
    .X(_07570_));
 sky130_fd_sc_hd__nor3_4 _24224_ (.A(_05302_),
    .B(_14316_),
    .C(_07479_),
    .Y(_07571_));
 sky130_fd_sc_hd__a41oi_4 _24225_ (.A1(_05403_),
    .A2(_05300_),
    .A3(_07570_),
    .A4(_07468_),
    .B1(_07571_),
    .Y(_07572_));
 sky130_fd_sc_hd__nor2_1 _24226_ (.A(_07483_),
    .B(_07490_),
    .Y(_07573_));
 sky130_fd_sc_hd__o21bai_4 _24227_ (.A1(_07480_),
    .A2(_07491_),
    .B1_N(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__clkbuf_4 _24228_ (.A(_07210_),
    .X(_07575_));
 sky130_fd_sc_hd__and2_2 _24229_ (.A(_14083_),
    .B(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__nand2_2 _24230_ (.A(_04905_),
    .B(_07477_),
    .Y(_07577_));
 sky130_fd_sc_hd__clkbuf_4 _24231_ (.A(_07484_),
    .X(_07578_));
 sky130_fd_sc_hd__nand2_2 _24232_ (.A(_04910_),
    .B(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__xnor2_4 _24233_ (.A(_07577_),
    .B(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__xor2_4 _24234_ (.A(_07576_),
    .B(_07580_),
    .X(_07581_));
 sky130_fd_sc_hd__nand3b_1 _24235_ (.A_N(_07487_),
    .B(_05420_),
    .C(_07034_),
    .Y(_07582_));
 sky130_fd_sc_hd__o31a_2 _24236_ (.A1(_05315_),
    .A2(_14298_),
    .A3(_07489_),
    .B1(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__buf_2 _24237_ (.A(\pcpi_mul.rs1[28] ),
    .X(_07584_));
 sky130_fd_sc_hd__clkbuf_4 _24238_ (.A(_07584_),
    .X(_07585_));
 sky130_fd_sc_hd__and2_2 _24239_ (.A(_05319_),
    .B(_07585_),
    .X(_07586_));
 sky130_fd_sc_hd__nand2_2 _24240_ (.A(_06445_),
    .B(_07038_),
    .Y(_07587_));
 sky130_fd_sc_hd__and2_1 _24241_ (.A(_05108_),
    .B(_07204_),
    .X(_07588_));
 sky130_fd_sc_hd__xor2_4 _24242_ (.A(_07587_),
    .B(_07588_),
    .X(_07589_));
 sky130_fd_sc_hd__xor2_4 _24243_ (.A(_07586_),
    .B(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__xnor2_4 _24244_ (.A(_07583_),
    .B(_07590_),
    .Y(_07591_));
 sky130_fd_sc_hd__xor2_4 _24245_ (.A(_07581_),
    .B(_07591_),
    .X(_07592_));
 sky130_fd_sc_hd__xnor2_4 _24246_ (.A(_07574_),
    .B(_07592_),
    .Y(_07593_));
 sky130_fd_sc_hd__xor2_4 _24247_ (.A(_07572_),
    .B(_07593_),
    .X(_07594_));
 sky130_fd_sc_hd__a21o_1 _24248_ (.A1(_07566_),
    .A2(_07567_),
    .B1(_07594_),
    .X(_07595_));
 sky130_fd_sc_hd__nand3_4 _24249_ (.A(_07566_),
    .B(_07594_),
    .C(_07567_),
    .Y(_07596_));
 sky130_fd_sc_hd__o21bai_2 _24250_ (.A1(_07431_),
    .A2(_07427_),
    .B1_N(_07428_),
    .Y(_07597_));
 sky130_fd_sc_hd__a21o_1 _24251_ (.A1(_07595_),
    .A2(_07596_),
    .B1(_07597_),
    .X(_07598_));
 sky130_fd_sc_hd__nand3_4 _24252_ (.A(_07595_),
    .B(_07597_),
    .C(_07596_),
    .Y(_07599_));
 sky130_fd_sc_hd__a21oi_1 _24253_ (.A1(_07466_),
    .A2(_07494_),
    .B1(_07463_),
    .Y(_07600_));
 sky130_vsdinv _24254_ (.A(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__a21o_1 _24255_ (.A1(_07598_),
    .A2(_07599_),
    .B1(_07601_),
    .X(_07602_));
 sky130_fd_sc_hd__nand3_4 _24256_ (.A(_07598_),
    .B(_07601_),
    .C(_07599_),
    .Y(_07603_));
 sky130_fd_sc_hd__nand2_2 _24257_ (.A(_07602_),
    .B(_07603_),
    .Y(_07604_));
 sky130_fd_sc_hd__nor2_1 _24258_ (.A(_07380_),
    .B(_07385_),
    .Y(_07605_));
 sky130_fd_sc_hd__o21ba_1 _24259_ (.A1(_07378_),
    .A2(_07386_),
    .B1_N(_07605_),
    .X(_07606_));
 sky130_fd_sc_hd__and2_2 _24260_ (.A(_06319_),
    .B(_05404_),
    .X(_07607_));
 sky130_fd_sc_hd__nand3_4 _24261_ (.A(_14009_),
    .B(_06737_),
    .C(_05427_),
    .Y(_07608_));
 sky130_fd_sc_hd__a22o_1 _24262_ (.A1(_06321_),
    .A2(_05105_),
    .B1(_06737_),
    .B2(_05236_),
    .X(_07609_));
 sky130_fd_sc_hd__o21ai_2 _24263_ (.A1(_06127_),
    .A2(_07608_),
    .B1(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__xnor2_2 _24264_ (.A(_07607_),
    .B(_07610_),
    .Y(_07611_));
 sky130_vsdinv _24265_ (.A(_07611_),
    .Y(_07612_));
 sky130_fd_sc_hd__a22o_1 _24266_ (.A1(_06744_),
    .A2(_05184_),
    .B1(_14001_),
    .B2(_05098_),
    .X(_07613_));
 sky130_fd_sc_hd__nand3_4 _24267_ (.A(_13997_),
    .B(\pcpi_mul.rs2[22] ),
    .C(_14426_),
    .Y(_07614_));
 sky130_fd_sc_hd__or2b_1 _24268_ (.A(_07614_),
    .B_N(_04983_),
    .X(_07615_));
 sky130_fd_sc_hd__o2bb2ai_1 _24269_ (.A1_N(_07613_),
    .A2_N(_07615_),
    .B1(_14004_),
    .B2(_14417_),
    .Y(_07616_));
 sky130_fd_sc_hd__o2111ai_4 _24270_ (.A1(_14421_),
    .A2(_07614_),
    .B1(_06470_),
    .C1(_05048_),
    .D1(_07613_),
    .Y(_07617_));
 sky130_fd_sc_hd__nand2_2 _24271_ (.A(_07616_),
    .B(_07617_),
    .Y(_07618_));
 sky130_fd_sc_hd__nand3b_1 _24272_ (.A_N(_07382_),
    .B(_07246_),
    .C(_04976_),
    .Y(_07619_));
 sky130_fd_sc_hd__o31a_1 _24273_ (.A1(_14005_),
    .A2(_14422_),
    .A3(_07384_),
    .B1(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__xnor2_1 _24274_ (.A(_07618_),
    .B(_07620_),
    .Y(_07621_));
 sky130_fd_sc_hd__xor2_1 _24275_ (.A(_07612_),
    .B(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__nor2_1 _24276_ (.A(_07362_),
    .B(_07367_),
    .Y(_07623_));
 sky130_fd_sc_hd__and2_2 _24277_ (.A(_07622_),
    .B(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__o21bai_4 _24278_ (.A1(_07367_),
    .A2(_07362_),
    .B1_N(_07622_),
    .Y(_07625_));
 sky130_fd_sc_hd__nor3b_4 _24279_ (.A(_07606_),
    .B(_07624_),
    .C_N(_07625_),
    .Y(_07626_));
 sky130_vsdinv _24280_ (.A(_07624_),
    .Y(_07627_));
 sky130_vsdinv _24281_ (.A(_07606_),
    .Y(_07628_));
 sky130_fd_sc_hd__a21oi_4 _24282_ (.A1(_07627_),
    .A2(_07625_),
    .B1(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__nor2_4 _24283_ (.A(_07361_),
    .B(_07368_),
    .Y(_07630_));
 sky130_fd_sc_hd__nand2_2 _24284_ (.A(_13976_),
    .B(_05533_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_2 _24285_ (.A(_07359_),
    .B(_04873_),
    .Y(_07632_));
 sky130_fd_sc_hd__xnor2_4 _24286_ (.A(_07631_),
    .B(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__o32a_4 _24287_ (.A1(_13993_),
    .A2(_05178_),
    .A3(_07366_),
    .B1(_14444_),
    .B2(_07263_),
    .X(_07634_));
 sky130_fd_sc_hd__nand2_2 _24288_ (.A(_06887_),
    .B(_04957_),
    .Y(_07635_));
 sky130_fd_sc_hd__or4_4 _24289_ (.A(_13984_),
    .B(_13988_),
    .C(_14437_),
    .D(_14442_),
    .X(_07636_));
 sky130_fd_sc_hd__a22o_1 _24290_ (.A1(_07261_),
    .A2(_04889_),
    .B1(_07265_),
    .B2(_05051_),
    .X(_07637_));
 sky130_fd_sc_hd__nand2_2 _24291_ (.A(_07636_),
    .B(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__xnor2_4 _24292_ (.A(_07635_),
    .B(_07638_),
    .Y(_07639_));
 sky130_fd_sc_hd__xnor2_4 _24293_ (.A(_07634_),
    .B(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__xor2_4 _24294_ (.A(_07633_),
    .B(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__xor2_1 _24295_ (.A(_07630_),
    .B(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__o21ba_1 _24296_ (.A1(_07626_),
    .A2(_07629_),
    .B1_N(_07642_),
    .X(_07643_));
 sky130_fd_sc_hd__nor3b_4 _24297_ (.A(_07626_),
    .B(_07629_),
    .C_N(_07642_),
    .Y(_07644_));
 sky130_vsdinv _24298_ (.A(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__nand3b_4 _24299_ (.A_N(_07643_),
    .B(_07645_),
    .C(_07391_),
    .Y(_07646_));
 sky130_fd_sc_hd__o2bb2ai_2 _24300_ (.A1_N(_07369_),
    .A2_N(_07389_),
    .B1(_07644_),
    .B2(_07643_),
    .Y(_07647_));
 sky130_fd_sc_hd__buf_2 _24301_ (.A(_14344_),
    .X(_07648_));
 sky130_fd_sc_hd__and2_2 _24302_ (.A(_05354_),
    .B(_07648_),
    .X(_07649_));
 sky130_fd_sc_hd__clkbuf_4 _24303_ (.A(_06028_),
    .X(_07650_));
 sky130_fd_sc_hd__nand3_4 _24304_ (.A(_05361_),
    .B(_05363_),
    .C(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__a22o_2 _24305_ (.A1(_05581_),
    .A2(_06029_),
    .B1(_06200_),
    .B2(_06154_),
    .X(_07652_));
 sky130_fd_sc_hd__o21ai_4 _24306_ (.A1(_14352_),
    .A2(_07651_),
    .B1(_07652_),
    .Y(_07653_));
 sky130_fd_sc_hd__xnor2_4 _24307_ (.A(_07649_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__buf_4 _24308_ (.A(_05635_),
    .X(_07655_));
 sky130_fd_sc_hd__nand3b_1 _24309_ (.A_N(_07402_),
    .B(_07655_),
    .C(_05512_),
    .Y(_07656_));
 sky130_fd_sc_hd__o31a_4 _24310_ (.A1(_14046_),
    .A2(_14371_),
    .A3(_07404_),
    .B1(_07656_),
    .X(_07657_));
 sky130_fd_sc_hd__and2_2 _24311_ (.A(_05440_),
    .B(_05776_),
    .X(_07658_));
 sky130_fd_sc_hd__nand2_2 _24312_ (.A(_06855_),
    .B(\pcpi_mul.rs1[15] ),
    .Y(_07659_));
 sky130_fd_sc_hd__and2_1 _24313_ (.A(_05634_),
    .B(\pcpi_mul.rs1[14] ),
    .X(_07660_));
 sky130_fd_sc_hd__xor2_4 _24314_ (.A(_07659_),
    .B(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__xor2_4 _24315_ (.A(_07658_),
    .B(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__xnor2_4 _24316_ (.A(_07657_),
    .B(_07662_),
    .Y(_07663_));
 sky130_fd_sc_hd__xnor2_4 _24317_ (.A(_07654_),
    .B(_07663_),
    .Y(_07664_));
 sky130_vsdinv _24318_ (.A(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__nor2_1 _24319_ (.A(_07414_),
    .B(_07419_),
    .Y(_07666_));
 sky130_fd_sc_hd__o21bai_2 _24320_ (.A1(_07412_),
    .A2(_07420_),
    .B1_N(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__buf_6 _24321_ (.A(_14389_),
    .X(_07668_));
 sky130_fd_sc_hd__nand3b_2 _24322_ (.A_N(_07416_),
    .B(_07295_),
    .C(_05406_),
    .Y(_07669_));
 sky130_fd_sc_hd__o31a_4 _24323_ (.A1(_14032_),
    .A2(_07668_),
    .A3(_07418_),
    .B1(_07669_),
    .X(_07670_));
 sky130_fd_sc_hd__a2bb2oi_4 _24324_ (.A1_N(_14411_),
    .A2_N(_07374_),
    .B1(_07373_),
    .B2(_07375_),
    .Y(_07671_));
 sky130_fd_sc_hd__and2_2 _24325_ (.A(\pcpi_mul.rs2[15] ),
    .B(_06040_),
    .X(_07672_));
 sky130_fd_sc_hd__nand2_2 _24326_ (.A(_06070_),
    .B(_14387_),
    .Y(_07673_));
 sky130_fd_sc_hd__and2_1 _24327_ (.A(_14022_),
    .B(\pcpi_mul.rs1[11] ),
    .X(_07674_));
 sky130_fd_sc_hd__xor2_4 _24328_ (.A(_07673_),
    .B(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__xor2_4 _24329_ (.A(_07672_),
    .B(_07675_),
    .X(_07676_));
 sky130_fd_sc_hd__xnor2_4 _24330_ (.A(_07671_),
    .B(_07676_),
    .Y(_07677_));
 sky130_fd_sc_hd__xor2_4 _24331_ (.A(_07670_),
    .B(_07677_),
    .X(_07678_));
 sky130_fd_sc_hd__xnor2_2 _24332_ (.A(_07667_),
    .B(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__nor2_4 _24333_ (.A(_07665_),
    .B(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__and2b_1 _24334_ (.A_N(_07372_),
    .B(_07387_),
    .X(_07681_));
 sky130_fd_sc_hd__o21ba_1 _24335_ (.A1(_07371_),
    .A2(_07388_),
    .B1_N(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__nand2_1 _24336_ (.A(_07679_),
    .B(_07665_),
    .Y(_07683_));
 sky130_fd_sc_hd__nor3b_4 _24337_ (.A(_07680_),
    .B(_07682_),
    .C_N(_07683_),
    .Y(_07684_));
 sky130_vsdinv _24338_ (.A(_07684_),
    .Y(_07685_));
 sky130_vsdinv _24339_ (.A(_07680_),
    .Y(_07686_));
 sky130_fd_sc_hd__a21bo_1 _24340_ (.A1(_07686_),
    .A2(_07683_),
    .B1_N(_07682_),
    .X(_07687_));
 sky130_fd_sc_hd__a21oi_1 _24341_ (.A1(_07421_),
    .A2(_07410_),
    .B1(_07423_),
    .Y(_07688_));
 sky130_vsdinv _24342_ (.A(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__a21o_1 _24343_ (.A1(_07685_),
    .A2(_07687_),
    .B1(_07689_),
    .X(_07690_));
 sky130_fd_sc_hd__nand3b_4 _24344_ (.A_N(_07684_),
    .B(_07689_),
    .C(_07687_),
    .Y(_07691_));
 sky130_fd_sc_hd__a22oi_4 _24345_ (.A1(_07646_),
    .A2(_07647_),
    .B1(_07690_),
    .B2(_07691_),
    .Y(_07692_));
 sky130_fd_sc_hd__nand2_2 _24346_ (.A(_07646_),
    .B(_07647_),
    .Y(_07693_));
 sky130_fd_sc_hd__nand2_2 _24347_ (.A(_07690_),
    .B(_07691_),
    .Y(_07694_));
 sky130_fd_sc_hd__nor2_4 _24348_ (.A(_07693_),
    .B(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__nor2_2 _24349_ (.A(_07692_),
    .B(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__o21ai_4 _24350_ (.A1(_07392_),
    .A2(_07437_),
    .B1(_07696_),
    .Y(_07697_));
 sky130_fd_sc_hd__o21ba_1 _24351_ (.A1(_07393_),
    .A2(_07435_),
    .B1_N(_07392_),
    .X(_07698_));
 sky130_fd_sc_hd__o21ai_4 _24352_ (.A1(_07692_),
    .A2(_07695_),
    .B1(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__nand3b_2 _24353_ (.A_N(_07604_),
    .B(_07697_),
    .C(_07699_),
    .Y(_07700_));
 sky130_fd_sc_hd__a211oi_4 _24354_ (.A1(_07321_),
    .A2(_07438_),
    .B1(_07436_),
    .C1(_07437_),
    .Y(_07701_));
 sky130_fd_sc_hd__a31o_1 _24355_ (.A1(_07504_),
    .A2(_07439_),
    .A3(_07503_),
    .B1(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__nand2_2 _24356_ (.A(_07697_),
    .B(_07699_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand2_1 _24357_ (.A(_07703_),
    .B(_07604_),
    .Y(_07704_));
 sky130_fd_sc_hd__nand3_4 _24358_ (.A(_07700_),
    .B(_07702_),
    .C(_07704_),
    .Y(_07705_));
 sky130_fd_sc_hd__a22oi_4 _24359_ (.A1(_07602_),
    .A2(_07603_),
    .B1(_07697_),
    .B2(_07699_),
    .Y(_07706_));
 sky130_fd_sc_hd__nor2_2 _24360_ (.A(_07604_),
    .B(_07703_),
    .Y(_07707_));
 sky130_fd_sc_hd__a31oi_4 _24361_ (.A1(_07504_),
    .A2(_07439_),
    .A3(_07503_),
    .B1(_07701_),
    .Y(_07708_));
 sky130_fd_sc_hd__o21ai_4 _24362_ (.A1(_07706_),
    .A2(_07707_),
    .B1(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__nor2_1 _24363_ (.A(_07470_),
    .B(_07493_),
    .Y(_07710_));
 sky130_fd_sc_hd__a21o_4 _24364_ (.A1(_07492_),
    .A2(_07472_),
    .B1(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__a21boi_4 _24365_ (.A1(_07503_),
    .A2(_07501_),
    .B1_N(_07711_),
    .Y(_07712_));
 sky130_fd_sc_hd__nand2_1 _24366_ (.A(_07503_),
    .B(_07501_),
    .Y(_07713_));
 sky130_fd_sc_hd__nor2_4 _24367_ (.A(_07711_),
    .B(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__o2bb2ai_4 _24368_ (.A1_N(_07705_),
    .A2_N(_07709_),
    .B1(_07712_),
    .B2(_07714_),
    .Y(_07715_));
 sky130_fd_sc_hd__nor2_2 _24369_ (.A(_07712_),
    .B(_07714_),
    .Y(_07716_));
 sky130_fd_sc_hd__nand3_4 _24370_ (.A(_07709_),
    .B(_07705_),
    .C(_07716_),
    .Y(_07717_));
 sky130_fd_sc_hd__nand2_1 _24371_ (.A(_07715_),
    .B(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__a21boi_2 _24372_ (.A1(_07510_),
    .A2(_07522_),
    .B1_N(_07517_),
    .Y(_07719_));
 sky130_fd_sc_hd__nand2_1 _24373_ (.A(_07718_),
    .B(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__nand2_2 _24374_ (.A(_07525_),
    .B(_07517_),
    .Y(_07721_));
 sky130_fd_sc_hd__nand3_4 _24375_ (.A(_07721_),
    .B(_07715_),
    .C(_07717_),
    .Y(_07722_));
 sky130_fd_sc_hd__a21boi_4 _24376_ (.A1(_07236_),
    .A2(_07232_),
    .B1_N(_07520_),
    .Y(_07723_));
 sky130_fd_sc_hd__a21oi_1 _24377_ (.A1(_07720_),
    .A2(_07722_),
    .B1(_07723_),
    .Y(_07724_));
 sky130_vsdinv _24378_ (.A(_07723_),
    .Y(_07725_));
 sky130_fd_sc_hd__a21oi_4 _24379_ (.A1(_07715_),
    .A2(_07717_),
    .B1(_07721_),
    .Y(_07726_));
 sky130_fd_sc_hd__nor2_2 _24380_ (.A(_07719_),
    .B(_07718_),
    .Y(_07727_));
 sky130_fd_sc_hd__nor3_2 _24381_ (.A(_07725_),
    .B(_07726_),
    .C(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__o21ai_2 _24382_ (.A1(_07530_),
    .A2(_07531_),
    .B1(_07528_),
    .Y(_07729_));
 sky130_fd_sc_hd__o21bai_1 _24383_ (.A1(_07724_),
    .A2(_07728_),
    .B1_N(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__o21bai_2 _24384_ (.A1(_07726_),
    .A2(_07727_),
    .B1_N(_07723_),
    .Y(_07731_));
 sky130_fd_sc_hd__nand3_2 _24385_ (.A(_07720_),
    .B(_07723_),
    .C(_07722_),
    .Y(_07732_));
 sky130_fd_sc_hd__nand3_4 _24386_ (.A(_07731_),
    .B(_07732_),
    .C(_07729_),
    .Y(_07733_));
 sky130_fd_sc_hd__and2_1 _24387_ (.A(_07730_),
    .B(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__nand2_1 _24388_ (.A(_07544_),
    .B(_07350_),
    .Y(_07735_));
 sky130_fd_sc_hd__nor2_1 _24389_ (.A(_07735_),
    .B(_07541_),
    .Y(_07736_));
 sky130_fd_sc_hd__nor2_1 _24390_ (.A(_06998_),
    .B(_07172_),
    .Y(_07737_));
 sky130_fd_sc_hd__nand2_2 _24391_ (.A(_07736_),
    .B(_07737_),
    .Y(_07738_));
 sky130_fd_sc_hd__a21oi_1 _24392_ (.A1(_07538_),
    .A2(_07539_),
    .B1(_07535_),
    .Y(_07739_));
 sky130_vsdinv _24393_ (.A(_07540_),
    .Y(_07740_));
 sky130_fd_sc_hd__nor2_1 _24394_ (.A(_07739_),
    .B(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__nand3_1 _24395_ (.A(_07741_),
    .B(_07352_),
    .C(_07356_),
    .Y(_07742_));
 sky130_fd_sc_hd__a21oi_1 _24396_ (.A1(_07351_),
    .A2(_07536_),
    .B1(_07740_),
    .Y(_07743_));
 sky130_fd_sc_hd__nand2_2 _24397_ (.A(_07742_),
    .B(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__o21bai_4 _24398_ (.A1(_07738_),
    .A2(_07006_),
    .B1_N(_07744_),
    .Y(_07745_));
 sky130_fd_sc_hd__xor2_1 _24399_ (.A(_07734_),
    .B(_07745_),
    .X(_02647_));
 sky130_fd_sc_hd__buf_4 _24400_ (.A(_06576_),
    .X(_07746_));
 sky130_fd_sc_hd__buf_6 _24401_ (.A(_07746_),
    .X(_07747_));
 sky130_fd_sc_hd__nand3b_1 _24402_ (.A_N(_07551_),
    .B(_05577_),
    .C(_07747_),
    .Y(_07748_));
 sky130_fd_sc_hd__o31a_4 _24403_ (.A1(_05576_),
    .A2(_14328_),
    .A3(_07553_),
    .B1(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__a2bb2oi_4 _24404_ (.A1_N(_14353_),
    .A2_N(_07651_),
    .B1(_07649_),
    .B2(_07652_),
    .Y(_07750_));
 sky130_fd_sc_hd__and2_2 _24405_ (.A(_05483_),
    .B(_07204_),
    .X(_07751_));
 sky130_fd_sc_hd__nand3_4 _24406_ (.A(_14062_),
    .B(_05163_),
    .C(_14331_),
    .Y(_07752_));
 sky130_fd_sc_hd__a22o_2 _24407_ (.A1(_05486_),
    .A2(\pcpi_mul.rs1[21] ),
    .B1(_14066_),
    .B2(\pcpi_mul.rs1[22] ),
    .X(_07753_));
 sky130_fd_sc_hd__o21ai_4 _24408_ (.A1(_14326_),
    .A2(_07752_),
    .B1(_07753_),
    .Y(_07754_));
 sky130_fd_sc_hd__xor2_4 _24409_ (.A(_07751_),
    .B(_07754_),
    .X(_07755_));
 sky130_fd_sc_hd__xnor2_4 _24410_ (.A(_07750_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__xor2_4 _24411_ (.A(_07749_),
    .B(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__or2b_1 _24412_ (.A(_07663_),
    .B_N(_07654_),
    .X(_07758_));
 sky130_fd_sc_hd__o21ai_4 _24413_ (.A1(_07662_),
    .A2(_07657_),
    .B1(_07758_),
    .Y(_07759_));
 sky130_fd_sc_hd__xnor2_2 _24414_ (.A(_07757_),
    .B(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__nor2_1 _24415_ (.A(_07549_),
    .B(_07554_),
    .Y(_07761_));
 sky130_fd_sc_hd__o21ba_4 _24416_ (.A1(_07547_),
    .A2(_07555_),
    .B1_N(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__nand2_2 _24417_ (.A(_07760_),
    .B(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__nor2_4 _24418_ (.A(_07762_),
    .B(_07760_),
    .Y(_07764_));
 sky130_vsdinv _24419_ (.A(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__a21o_1 _24420_ (.A1(_07558_),
    .A2(_07556_),
    .B1(_07563_),
    .X(_07766_));
 sky130_fd_sc_hd__a21o_2 _24421_ (.A1(_07763_),
    .A2(_07765_),
    .B1(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__nand3_4 _24422_ (.A(_07766_),
    .B(_07765_),
    .C(_07763_),
    .Y(_07768_));
 sky130_fd_sc_hd__buf_4 _24423_ (.A(_07578_),
    .X(_07769_));
 sky130_fd_sc_hd__buf_4 _24424_ (.A(_07769_),
    .X(_07770_));
 sky130_fd_sc_hd__nor3_4 _24425_ (.A(_14087_),
    .B(_14311_),
    .C(_07580_),
    .Y(_07771_));
 sky130_fd_sc_hd__a41oi_4 _24426_ (.A1(_05403_),
    .A2(_05899_),
    .A3(_07770_),
    .A4(_07570_),
    .B1(_07771_),
    .Y(_07772_));
 sky130_fd_sc_hd__nor2_1 _24427_ (.A(_07583_),
    .B(_07590_),
    .Y(_07773_));
 sky130_fd_sc_hd__o21bai_4 _24428_ (.A1(_07581_),
    .A2(_07591_),
    .B1_N(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__buf_2 _24429_ (.A(_07568_),
    .X(_07775_));
 sky130_fd_sc_hd__and2_2 _24430_ (.A(_14083_),
    .B(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__nand2_2 _24431_ (.A(_04936_),
    .B(_07578_),
    .Y(_07777_));
 sky130_fd_sc_hd__buf_2 _24432_ (.A(_07584_),
    .X(_07778_));
 sky130_fd_sc_hd__nand2_2 _24433_ (.A(_04938_),
    .B(_07778_),
    .Y(_07779_));
 sky130_fd_sc_hd__xnor2_4 _24434_ (.A(_07777_),
    .B(_07779_),
    .Y(_07780_));
 sky130_fd_sc_hd__xor2_4 _24435_ (.A(_07776_),
    .B(_07780_),
    .X(_07781_));
 sky130_fd_sc_hd__nand3b_1 _24436_ (.A_N(_07587_),
    .B(_06159_),
    .C(_07206_),
    .Y(_07782_));
 sky130_fd_sc_hd__o31a_2 _24437_ (.A1(_14097_),
    .A2(_14292_),
    .A3(_07589_),
    .B1(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__buf_2 _24438_ (.A(\pcpi_mul.rs1[29] ),
    .X(_07784_));
 sky130_fd_sc_hd__and2_2 _24439_ (.A(_04955_),
    .B(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__buf_2 _24440_ (.A(\pcpi_mul.rs1[25] ),
    .X(_07786_));
 sky130_fd_sc_hd__nand2_4 _24441_ (.A(_06445_),
    .B(_07786_),
    .Y(_07787_));
 sky130_fd_sc_hd__and2_1 _24442_ (.A(_05108_),
    .B(_06956_),
    .X(_07788_));
 sky130_fd_sc_hd__xor2_4 _24443_ (.A(_07787_),
    .B(_07788_),
    .X(_07789_));
 sky130_fd_sc_hd__xor2_4 _24444_ (.A(_07785_),
    .B(_07789_),
    .X(_07790_));
 sky130_fd_sc_hd__xnor2_4 _24445_ (.A(_07783_),
    .B(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__xor2_4 _24446_ (.A(_07781_),
    .B(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__xnor2_4 _24447_ (.A(_07774_),
    .B(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__xor2_4 _24448_ (.A(_07772_),
    .B(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__a21o_1 _24449_ (.A1(_07767_),
    .A2(_07768_),
    .B1(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__nand3_4 _24450_ (.A(_07767_),
    .B(_07794_),
    .C(_07768_),
    .Y(_07796_));
 sky130_fd_sc_hd__a21o_1 _24451_ (.A1(_07687_),
    .A2(_07689_),
    .B1(_07684_),
    .X(_07797_));
 sky130_fd_sc_hd__a21o_2 _24452_ (.A1(_07795_),
    .A2(_07796_),
    .B1(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__nand3_4 _24453_ (.A(_07795_),
    .B(_07797_),
    .C(_07796_),
    .Y(_07799_));
 sky130_fd_sc_hd__a21boi_1 _24454_ (.A1(_07566_),
    .A2(_07594_),
    .B1_N(_07567_),
    .Y(_07800_));
 sky130_vsdinv _24455_ (.A(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__a21o_1 _24456_ (.A1(_07798_),
    .A2(_07799_),
    .B1(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__nand3_4 _24457_ (.A(_07798_),
    .B(_07801_),
    .C(_07799_),
    .Y(_07803_));
 sky130_fd_sc_hd__and2_2 _24458_ (.A(_05354_),
    .B(_06576_),
    .X(_07804_));
 sky130_fd_sc_hd__nand3_4 _24459_ (.A(_05879_),
    .B(_06200_),
    .C(_06037_),
    .Y(_07805_));
 sky130_fd_sc_hd__a22o_2 _24460_ (.A1(_05358_),
    .A2(_06287_),
    .B1(_06202_),
    .B2(_07648_),
    .X(_07806_));
 sky130_fd_sc_hd__o21ai_4 _24461_ (.A1(_06293_),
    .A2(_07805_),
    .B1(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__xnor2_4 _24462_ (.A(_07804_),
    .B(_07807_),
    .Y(_07808_));
 sky130_fd_sc_hd__a22o_1 _24463_ (.A1(_05730_),
    .A2(\pcpi_mul.rs1[15] ),
    .B1(_06855_),
    .B2(_06017_),
    .X(_07809_));
 sky130_fd_sc_hd__nand3_4 _24464_ (.A(_05954_),
    .B(_14040_),
    .C(\pcpi_mul.rs1[15] ),
    .Y(_07810_));
 sky130_fd_sc_hd__or2b_1 _24465_ (.A(_07810_),
    .B_N(_05776_),
    .X(_07811_));
 sky130_fd_sc_hd__o2bb2ai_1 _24466_ (.A1_N(_07809_),
    .A2_N(_07811_),
    .B1(_06206_),
    .B2(_14358_),
    .Y(_07812_));
 sky130_fd_sc_hd__o2111ai_4 _24467_ (.A1(_14364_),
    .A2(_07810_),
    .B1(_05728_),
    .C1(_05912_),
    .D1(_07809_),
    .Y(_07813_));
 sky130_fd_sc_hd__and2_2 _24468_ (.A(_07812_),
    .B(_07813_),
    .X(_07814_));
 sky130_fd_sc_hd__nand3b_1 _24469_ (.A_N(_07659_),
    .B(_07281_),
    .C(_05610_),
    .Y(_07815_));
 sky130_fd_sc_hd__o31a_2 _24470_ (.A1(_06207_),
    .A2(_14365_),
    .A3(_07661_),
    .B1(_07815_),
    .X(_07816_));
 sky130_fd_sc_hd__xor2_4 _24471_ (.A(_07814_),
    .B(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__xnor2_4 _24472_ (.A(_07808_),
    .B(_07817_),
    .Y(_07818_));
 sky130_vsdinv _24473_ (.A(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__buf_6 _24474_ (.A(_06067_),
    .X(_07820_));
 sky130_fd_sc_hd__nand3b_2 _24475_ (.A_N(_07673_),
    .B(_07820_),
    .C(_05498_),
    .Y(_07821_));
 sky130_fd_sc_hd__o31a_4 _24476_ (.A1(_14032_),
    .A2(_06409_),
    .A3(_07675_),
    .B1(_07821_),
    .X(_07822_));
 sky130_fd_sc_hd__a2bb2oi_4 _24477_ (.A1_N(_06127_),
    .A2_N(_07608_),
    .B1(_07607_),
    .B2(_07609_),
    .Y(_07823_));
 sky130_fd_sc_hd__a22o_1 _24478_ (.A1(_06348_),
    .A2(_05917_),
    .B1(_06351_),
    .B2(_06040_),
    .X(_07824_));
 sky130_fd_sc_hd__nand3_4 _24479_ (.A(_06485_),
    .B(_14026_),
    .C(_14387_),
    .Y(_07825_));
 sky130_fd_sc_hd__or2b_1 _24480_ (.A(_07825_),
    .B_N(_05915_),
    .X(_07826_));
 sky130_fd_sc_hd__o2bb2ai_1 _24481_ (.A1_N(_07824_),
    .A2_N(_07826_),
    .B1(_14031_),
    .B2(_14378_),
    .Y(_07827_));
 sky130_fd_sc_hd__o2111ai_4 _24482_ (.A1(_14383_),
    .A2(_07825_),
    .B1(_06489_),
    .C1(_05610_),
    .D1(_07824_),
    .Y(_07828_));
 sky130_fd_sc_hd__nand2_4 _24483_ (.A(_07827_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__xnor2_4 _24484_ (.A(_07823_),
    .B(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__xor2_4 _24485_ (.A(_07822_),
    .B(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__nor2_1 _24486_ (.A(_07671_),
    .B(_07676_),
    .Y(_07832_));
 sky130_fd_sc_hd__o21bai_2 _24487_ (.A1(_07670_),
    .A2(_07677_),
    .B1_N(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__xnor2_2 _24488_ (.A(_07831_),
    .B(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__nor2_4 _24489_ (.A(_07819_),
    .B(_07834_),
    .Y(_07835_));
 sky130_fd_sc_hd__a21oi_4 _24490_ (.A1(_07625_),
    .A2(_07628_),
    .B1(_07624_),
    .Y(_07836_));
 sky130_fd_sc_hd__nand2_1 _24491_ (.A(_07834_),
    .B(_07819_),
    .Y(_07837_));
 sky130_fd_sc_hd__nor3b_4 _24492_ (.A(_07835_),
    .B(_07836_),
    .C_N(_07837_),
    .Y(_07838_));
 sky130_vsdinv _24493_ (.A(_07838_),
    .Y(_07839_));
 sky130_vsdinv _24494_ (.A(_07835_),
    .Y(_07840_));
 sky130_fd_sc_hd__a21bo_1 _24495_ (.A1(_07840_),
    .A2(_07837_),
    .B1_N(_07836_),
    .X(_07841_));
 sky130_fd_sc_hd__a21oi_1 _24496_ (.A1(_07678_),
    .A2(_07667_),
    .B1(_07680_),
    .Y(_07842_));
 sky130_vsdinv _24497_ (.A(_07842_),
    .Y(_07843_));
 sky130_fd_sc_hd__a21o_1 _24498_ (.A1(_07839_),
    .A2(_07841_),
    .B1(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__nand3b_1 _24499_ (.A_N(_07838_),
    .B(_07843_),
    .C(_07841_),
    .Y(_07845_));
 sky130_fd_sc_hd__nand2_2 _24500_ (.A(_07844_),
    .B(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__nor2_1 _24501_ (.A(_07618_),
    .B(_07620_),
    .Y(_07847_));
 sky130_fd_sc_hd__o21ba_1 _24502_ (.A1(_07612_),
    .A2(_07621_),
    .B1_N(_07847_),
    .X(_07848_));
 sky130_fd_sc_hd__and2_2 _24503_ (.A(_06319_),
    .B(_05413_),
    .X(_07849_));
 sky130_fd_sc_hd__nand3_4 _24504_ (.A(_14009_),
    .B(_14014_),
    .C(_05308_),
    .Y(_07850_));
 sky130_fd_sc_hd__a22o_1 _24505_ (.A1(_06321_),
    .A2(_05181_),
    .B1(_06737_),
    .B2(_05404_),
    .X(_07851_));
 sky130_fd_sc_hd__o21ai_2 _24506_ (.A1(_14400_),
    .A2(_07850_),
    .B1(_07851_),
    .Y(_07852_));
 sky130_fd_sc_hd__xnor2_2 _24507_ (.A(_07849_),
    .B(_07852_),
    .Y(_07853_));
 sky130_vsdinv _24508_ (.A(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__o21a_1 _24509_ (.A1(_14422_),
    .A2(_07614_),
    .B1(_07617_),
    .X(_07855_));
 sky130_fd_sc_hd__a22o_1 _24510_ (.A1(_13998_),
    .A2(_04983_),
    .B1(_06646_),
    .B2(_05429_),
    .X(_07856_));
 sky130_fd_sc_hd__nand3_4 _24511_ (.A(_13997_),
    .B(_14001_),
    .C(_05090_),
    .Y(_07857_));
 sky130_fd_sc_hd__or2b_1 _24512_ (.A(_07857_),
    .B_N(_05429_),
    .X(_07858_));
 sky130_fd_sc_hd__o2bb2ai_1 _24513_ (.A1_N(_07856_),
    .A2_N(_07858_),
    .B1(_14005_),
    .B2(_05998_),
    .Y(_07859_));
 sky130_fd_sc_hd__o2111ai_4 _24514_ (.A1(_14417_),
    .A2(_07857_),
    .B1(_06470_),
    .C1(_05228_),
    .D1(_07856_),
    .Y(_07860_));
 sky130_fd_sc_hd__nand2_2 _24515_ (.A(_07859_),
    .B(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__xnor2_1 _24516_ (.A(_07855_),
    .B(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__xor2_1 _24517_ (.A(_07854_),
    .B(_07862_),
    .X(_07863_));
 sky130_fd_sc_hd__nor2_1 _24518_ (.A(_07634_),
    .B(_07639_),
    .Y(_07864_));
 sky130_fd_sc_hd__and2_2 _24519_ (.A(_07863_),
    .B(_07864_),
    .X(_07865_));
 sky130_fd_sc_hd__o21bai_4 _24520_ (.A1(_07634_),
    .A2(_07639_),
    .B1_N(_07863_),
    .Y(_07866_));
 sky130_fd_sc_hd__nor3b_4 _24521_ (.A(_07848_),
    .B(_07865_),
    .C_N(_07866_),
    .Y(_07867_));
 sky130_vsdinv _24522_ (.A(_07865_),
    .Y(_07868_));
 sky130_vsdinv _24523_ (.A(_07848_),
    .Y(_07869_));
 sky130_fd_sc_hd__a21oi_4 _24524_ (.A1(_07868_),
    .A2(_07866_),
    .B1(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__nor2_1 _24525_ (.A(_07633_),
    .B(_07640_),
    .Y(_07871_));
 sky130_vsdinv _24526_ (.A(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__buf_4 _24527_ (.A(\pcpi_mul.rs2[27] ),
    .X(_07873_));
 sky130_fd_sc_hd__and2_1 _24528_ (.A(_07873_),
    .B(_04891_),
    .X(_07874_));
 sky130_fd_sc_hd__nand2_2 _24529_ (.A(\pcpi_mul.rs2[28] ),
    .B(_04986_),
    .Y(_07875_));
 sky130_fd_sc_hd__nand2_1 _24530_ (.A(\pcpi_mul.rs2[29] ),
    .B(_04716_),
    .Y(_07876_));
 sky130_fd_sc_hd__xnor2_2 _24531_ (.A(_07875_),
    .B(_07876_),
    .Y(_07877_));
 sky130_fd_sc_hd__xnor2_2 _24532_ (.A(_07874_),
    .B(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__o21a_2 _24533_ (.A1(_07635_),
    .A2(_07638_),
    .B1(_07636_),
    .X(_07879_));
 sky130_fd_sc_hd__nand3b_4 _24534_ (.A_N(_07631_),
    .B(\pcpi_mul.rs2[27] ),
    .C(_04872_),
    .Y(_07880_));
 sky130_fd_sc_hd__a22o_1 _24535_ (.A1(_07261_),
    .A2(_04897_),
    .B1(_07101_),
    .B2(_14432_),
    .X(_07881_));
 sky130_fd_sc_hd__nand3_4 _24536_ (.A(\pcpi_mul.rs2[26] ),
    .B(\pcpi_mul.rs2[25] ),
    .C(_04948_),
    .Y(_07882_));
 sky130_fd_sc_hd__or2b_1 _24537_ (.A(_07882_),
    .B_N(_04956_),
    .X(_07883_));
 sky130_fd_sc_hd__o2bb2ai_2 _24538_ (.A1_N(_07881_),
    .A2_N(_07883_),
    .B1(_13993_),
    .B2(_14428_),
    .Y(_07884_));
 sky130_fd_sc_hd__o2111ai_4 _24539_ (.A1(_14433_),
    .A2(_07882_),
    .B1(\pcpi_mul.rs2[24] ),
    .C1(_04978_),
    .D1(_07881_),
    .Y(_07885_));
 sky130_fd_sc_hd__nand2_2 _24540_ (.A(_07884_),
    .B(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__xnor2_4 _24541_ (.A(_07880_),
    .B(_07886_),
    .Y(_07887_));
 sky130_fd_sc_hd__xor2_2 _24542_ (.A(_07879_),
    .B(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__xnor2_1 _24543_ (.A(_07878_),
    .B(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__nor2_2 _24544_ (.A(_07872_),
    .B(_07889_),
    .Y(_07890_));
 sky130_fd_sc_hd__o21a_1 _24545_ (.A1(_07633_),
    .A2(_07640_),
    .B1(_07889_),
    .X(_07891_));
 sky130_fd_sc_hd__o22a_1 _24546_ (.A1(_07867_),
    .A2(_07870_),
    .B1(_07890_),
    .B2(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__nor2_1 _24547_ (.A(_07890_),
    .B(_07891_),
    .Y(_07893_));
 sky130_fd_sc_hd__nor3b_4 _24548_ (.A(_07867_),
    .B(_07870_),
    .C_N(_07893_),
    .Y(_07894_));
 sky130_fd_sc_hd__nor2_4 _24549_ (.A(_07892_),
    .B(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__a211oi_4 _24550_ (.A1(_07630_),
    .A2(_07641_),
    .B1(_07644_),
    .C1(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__a21o_1 _24551_ (.A1(_07630_),
    .A2(_07641_),
    .B1(_07644_),
    .X(_07897_));
 sky130_fd_sc_hd__nand2_1 _24552_ (.A(_07897_),
    .B(_07895_),
    .Y(_07898_));
 sky130_fd_sc_hd__nor3b_4 _24553_ (.A(_07846_),
    .B(_07896_),
    .C_N(_07898_),
    .Y(_07899_));
 sky130_vsdinv _24554_ (.A(_07898_),
    .Y(_07900_));
 sky130_fd_sc_hd__o21a_1 _24555_ (.A1(_07896_),
    .A2(_07900_),
    .B1(_07846_),
    .X(_07901_));
 sky130_fd_sc_hd__o21ai_2 _24556_ (.A1(_07693_),
    .A2(_07694_),
    .B1(_07646_),
    .Y(_07902_));
 sky130_fd_sc_hd__o21bai_4 _24557_ (.A1(_07899_),
    .A2(_07901_),
    .B1_N(_07902_),
    .Y(_07903_));
 sky130_vsdinv _24558_ (.A(_07899_),
    .Y(_07904_));
 sky130_fd_sc_hd__nand3b_4 _24559_ (.A_N(_07901_),
    .B(_07904_),
    .C(_07902_),
    .Y(_07905_));
 sky130_fd_sc_hd__a22oi_4 _24560_ (.A1(_07802_),
    .A2(_07803_),
    .B1(_07903_),
    .B2(_07905_),
    .Y(_07906_));
 sky130_fd_sc_hd__nand2_2 _24561_ (.A(_07802_),
    .B(_07803_),
    .Y(_07907_));
 sky130_fd_sc_hd__nand2_1 _24562_ (.A(_07903_),
    .B(_07905_),
    .Y(_07908_));
 sky130_fd_sc_hd__nor2_2 _24563_ (.A(_07907_),
    .B(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__o21a_1 _24564_ (.A1(_07604_),
    .A2(_07703_),
    .B1(_07697_),
    .X(_07910_));
 sky130_fd_sc_hd__o21ai_4 _24565_ (.A1(_07906_),
    .A2(_07909_),
    .B1(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__o21ai_2 _24566_ (.A1(_07604_),
    .A2(_07703_),
    .B1(_07697_),
    .Y(_07912_));
 sky130_fd_sc_hd__nand3b_4 _24567_ (.A_N(_07907_),
    .B(_07905_),
    .C(_07903_),
    .Y(_07913_));
 sky130_fd_sc_hd__nand2_2 _24568_ (.A(_07908_),
    .B(_07907_),
    .Y(_07914_));
 sky130_fd_sc_hd__nand3_4 _24569_ (.A(_07912_),
    .B(_07913_),
    .C(_07914_),
    .Y(_07915_));
 sky130_fd_sc_hd__nor2_2 _24570_ (.A(_07572_),
    .B(_07593_),
    .Y(_07916_));
 sky130_fd_sc_hd__a21oi_4 _24571_ (.A1(_07592_),
    .A2(_07574_),
    .B1(_07916_),
    .Y(_07917_));
 sky130_fd_sc_hd__a21oi_4 _24572_ (.A1(_07603_),
    .A2(_07599_),
    .B1(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__and3_2 _24573_ (.A(_07603_),
    .B(_07599_),
    .C(_07917_),
    .X(_07919_));
 sky130_fd_sc_hd__nor2_4 _24574_ (.A(_07918_),
    .B(_07919_),
    .Y(_07920_));
 sky130_fd_sc_hd__a21oi_1 _24575_ (.A1(_07911_),
    .A2(_07915_),
    .B1(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__nand3_4 _24576_ (.A(_07911_),
    .B(_07915_),
    .C(_07920_),
    .Y(_07922_));
 sky130_vsdinv _24577_ (.A(_07922_),
    .Y(_07923_));
 sky130_vsdinv _24578_ (.A(_07716_),
    .Y(_07924_));
 sky130_fd_sc_hd__o21a_1 _24579_ (.A1(_07706_),
    .A2(_07707_),
    .B1(_07708_),
    .X(_07925_));
 sky130_fd_sc_hd__o21ai_4 _24580_ (.A1(_07924_),
    .A2(_07925_),
    .B1(_07705_),
    .Y(_07926_));
 sky130_fd_sc_hd__o21bai_2 _24581_ (.A1(_07921_),
    .A2(_07923_),
    .B1_N(_07926_),
    .Y(_07927_));
 sky130_fd_sc_hd__clkbuf_4 _24582_ (.A(_07918_),
    .X(_07928_));
 sky130_fd_sc_hd__o2bb2ai_4 _24583_ (.A1_N(_07915_),
    .A2_N(_07911_),
    .B1(_07928_),
    .B2(_07919_),
    .Y(_07929_));
 sky130_fd_sc_hd__nand3_4 _24584_ (.A(_07929_),
    .B(_07926_),
    .C(_07922_),
    .Y(_07930_));
 sky130_fd_sc_hd__a21oi_2 _24585_ (.A1(_07927_),
    .A2(_07930_),
    .B1(_07712_),
    .Y(_07931_));
 sky130_fd_sc_hd__nand3_4 _24586_ (.A(_07927_),
    .B(_07930_),
    .C(_07712_),
    .Y(_07932_));
 sky130_vsdinv _24587_ (.A(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__o21ai_4 _24588_ (.A1(_07725_),
    .A2(_07726_),
    .B1(_07722_),
    .Y(_07934_));
 sky130_fd_sc_hd__o21bai_1 _24589_ (.A1(_07931_),
    .A2(_07933_),
    .B1_N(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__a21oi_4 _24590_ (.A1(_07929_),
    .A2(_07922_),
    .B1(_07926_),
    .Y(_07936_));
 sky130_vsdinv _24591_ (.A(_07930_),
    .Y(_07937_));
 sky130_fd_sc_hd__o21bai_4 _24592_ (.A1(_07936_),
    .A2(_07937_),
    .B1_N(_07712_),
    .Y(_07938_));
 sky130_fd_sc_hd__nand3_4 _24593_ (.A(_07938_),
    .B(_07934_),
    .C(_07932_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand2_2 _24594_ (.A(_07935_),
    .B(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__a21boi_1 _24595_ (.A1(_07745_),
    .A2(_07730_),
    .B1_N(_07733_),
    .Y(_07941_));
 sky130_fd_sc_hd__xor2_1 _24596_ (.A(_07940_),
    .B(_07941_),
    .X(_02648_));
 sky130_fd_sc_hd__o21a_1 _24597_ (.A1(_07846_),
    .A2(_07896_),
    .B1(_07898_),
    .X(_07942_));
 sky130_vsdinv _24598_ (.A(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__nand2_2 _24599_ (.A(_07888_),
    .B(_07878_),
    .Y(_07944_));
 sky130_fd_sc_hd__buf_4 _24600_ (.A(\pcpi_mul.rs2[30] ),
    .X(_07945_));
 sky130_fd_sc_hd__buf_4 _24601_ (.A(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__and2_2 _24602_ (.A(_07946_),
    .B(_04718_),
    .X(_07947_));
 sky130_fd_sc_hd__nand2_2 _24603_ (.A(_07358_),
    .B(_04974_),
    .Y(_07948_));
 sky130_fd_sc_hd__nand3b_2 _24604_ (.A_N(_07875_),
    .B(_13971_),
    .C(_04890_),
    .Y(_07949_));
 sky130_fd_sc_hd__a22o_1 _24605_ (.A1(\pcpi_mul.rs2[29] ),
    .A2(_04906_),
    .B1(_13976_),
    .B2(_04968_),
    .X(_07950_));
 sky130_fd_sc_hd__nand2_2 _24606_ (.A(_07949_),
    .B(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__xnor2_4 _24607_ (.A(_07948_),
    .B(_07951_),
    .Y(_07952_));
 sky130_fd_sc_hd__xnor2_4 _24608_ (.A(_07947_),
    .B(_07952_),
    .Y(_07953_));
 sky130_fd_sc_hd__o21a_2 _24609_ (.A1(_14435_),
    .A2(_07882_),
    .B1(_07885_),
    .X(_07954_));
 sky130_fd_sc_hd__a22o_1 _24610_ (.A1(_07261_),
    .A2(_05111_),
    .B1(_07101_),
    .B2(_04960_),
    .X(_07955_));
 sky130_fd_sc_hd__nand3_4 _24611_ (.A(_07261_),
    .B(_07101_),
    .C(_14432_),
    .Y(_07956_));
 sky130_fd_sc_hd__or2b_1 _24612_ (.A(_07956_),
    .B_N(_05959_),
    .X(_07957_));
 sky130_fd_sc_hd__o2bb2ai_1 _24613_ (.A1_N(_07955_),
    .A2_N(_07957_),
    .B1(_13993_),
    .B2(_14422_),
    .Y(_07958_));
 sky130_fd_sc_hd__o2111ai_4 _24614_ (.A1(_14427_),
    .A2(_07956_),
    .B1(_06887_),
    .C1(_05091_),
    .D1(_07955_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand2_4 _24615_ (.A(_07958_),
    .B(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__clkbuf_4 _24616_ (.A(\pcpi_mul.rs2[29] ),
    .X(_07961_));
 sky130_fd_sc_hd__nand3b_1 _24617_ (.A_N(_07875_),
    .B(_07961_),
    .C(_04717_),
    .Y(_07962_));
 sky130_fd_sc_hd__o31a_2 _24618_ (.A1(_13982_),
    .A2(_14443_),
    .A3(_07877_),
    .B1(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__xnor2_4 _24619_ (.A(_07960_),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__xor2_4 _24620_ (.A(_07954_),
    .B(_07964_),
    .X(_07965_));
 sky130_fd_sc_hd__xnor2_2 _24621_ (.A(_07953_),
    .B(_07965_),
    .Y(_07966_));
 sky130_fd_sc_hd__nor2_4 _24622_ (.A(_07944_),
    .B(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__and2_1 _24623_ (.A(_07966_),
    .B(_07944_),
    .X(_07968_));
 sky130_fd_sc_hd__nor2_1 _24624_ (.A(_07855_),
    .B(_07861_),
    .Y(_07969_));
 sky130_fd_sc_hd__o21ba_2 _24625_ (.A1(_07854_),
    .A2(_07862_),
    .B1_N(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__nand3b_2 _24626_ (.A_N(_07880_),
    .B(_07884_),
    .C(_07885_),
    .Y(_07971_));
 sky130_fd_sc_hd__o21ai_4 _24627_ (.A1(_07879_),
    .A2(_07887_),
    .B1(_07971_),
    .Y(_07972_));
 sky130_fd_sc_hd__and2_2 _24628_ (.A(_06319_),
    .B(_05423_),
    .X(_07973_));
 sky130_fd_sc_hd__nand3_4 _24629_ (.A(_14010_),
    .B(_06185_),
    .C(_05405_),
    .Y(_07974_));
 sky130_fd_sc_hd__a22o_2 _24630_ (.A1(_06322_),
    .A2(_05241_),
    .B1(_14014_),
    .B2(_05413_),
    .X(_07975_));
 sky130_fd_sc_hd__o21ai_4 _24631_ (.A1(_05418_),
    .A2(_07974_),
    .B1(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__xor2_4 _24632_ (.A(_07973_),
    .B(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__o21a_2 _24633_ (.A1(_05115_),
    .A2(_07857_),
    .B1(_07860_),
    .X(_07978_));
 sky130_fd_sc_hd__buf_2 _24634_ (.A(\pcpi_mul.rs2[22] ),
    .X(_07979_));
 sky130_fd_sc_hd__a22o_1 _24635_ (.A1(_13998_),
    .A2(_05047_),
    .B1(_07979_),
    .B2(_05105_),
    .X(_07980_));
 sky130_fd_sc_hd__nand3_4 _24636_ (.A(_13998_),
    .B(_06646_),
    .C(_05047_),
    .Y(_07981_));
 sky130_fd_sc_hd__or2b_1 _24637_ (.A(_07981_),
    .B_N(_05106_),
    .X(_07982_));
 sky130_fd_sc_hd__o2bb2ai_1 _24638_ (.A1_N(_07980_),
    .A2_N(_07982_),
    .B1(_14005_),
    .B2(_14405_),
    .Y(_07983_));
 sky130_fd_sc_hd__o2111ai_4 _24639_ (.A1(_05998_),
    .A2(_07981_),
    .B1(_06470_),
    .C1(_05237_),
    .D1(_07980_),
    .Y(_07984_));
 sky130_fd_sc_hd__nand2_4 _24640_ (.A(_07983_),
    .B(_07984_),
    .Y(_07985_));
 sky130_fd_sc_hd__xnor2_4 _24641_ (.A(_07978_),
    .B(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__xor2_4 _24642_ (.A(_07977_),
    .B(_07986_),
    .X(_07987_));
 sky130_fd_sc_hd__xnor2_4 _24643_ (.A(_07972_),
    .B(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__xor2_4 _24644_ (.A(_07970_),
    .B(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__nor3b_4 _24645_ (.A(_07967_),
    .B(_07968_),
    .C_N(_07989_),
    .Y(_07990_));
 sky130_fd_sc_hd__o21ba_1 _24646_ (.A1(_07967_),
    .A2(_07968_),
    .B1_N(_07989_),
    .X(_07991_));
 sky130_fd_sc_hd__nor2_2 _24647_ (.A(_07890_),
    .B(_07894_),
    .Y(_07992_));
 sky130_fd_sc_hd__or3_4 _24648_ (.A(_07990_),
    .B(_07991_),
    .C(_07992_),
    .X(_07993_));
 sky130_fd_sc_hd__o21ai_2 _24649_ (.A1(_07991_),
    .A2(_07990_),
    .B1(_07992_),
    .Y(_07994_));
 sky130_fd_sc_hd__nand2_1 _24650_ (.A(_07993_),
    .B(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__a21oi_1 _24651_ (.A1(_07831_),
    .A2(_07833_),
    .B1(_07835_),
    .Y(_07996_));
 sky130_vsdinv _24652_ (.A(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__a21oi_4 _24653_ (.A1(_07866_),
    .A2(_07869_),
    .B1(_07865_),
    .Y(_07998_));
 sky130_fd_sc_hd__and2_2 _24654_ (.A(_05354_),
    .B(_07048_),
    .X(_07999_));
 sky130_fd_sc_hd__nand3_4 _24655_ (.A(_05879_),
    .B(_06200_),
    .C(_06583_),
    .Y(_08000_));
 sky130_fd_sc_hd__a22o_2 _24656_ (.A1(_05581_),
    .A2(_07648_),
    .B1(_06202_),
    .B2(_06296_),
    .X(_08001_));
 sky130_fd_sc_hd__o21ai_4 _24657_ (.A1(_14339_),
    .A2(_08000_),
    .B1(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__xnor2_4 _24658_ (.A(_07999_),
    .B(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__o21a_2 _24659_ (.A1(_14365_),
    .A2(_07810_),
    .B1(_07813_),
    .X(_08004_));
 sky130_fd_sc_hd__a22o_1 _24660_ (.A1(_14036_),
    .A2(_06017_),
    .B1(_05732_),
    .B2(_14357_),
    .X(_08005_));
 sky130_fd_sc_hd__nand3_4 _24661_ (.A(_05954_),
    .B(_06855_),
    .C(\pcpi_mul.rs1[16] ),
    .Y(_08006_));
 sky130_fd_sc_hd__or2b_1 _24662_ (.A(_08006_),
    .B_N(_06028_),
    .X(_08007_));
 sky130_fd_sc_hd__o2bb2ai_1 _24663_ (.A1_N(_08005_),
    .A2_N(_08007_),
    .B1(_14046_),
    .B2(_14351_),
    .Y(_08008_));
 sky130_fd_sc_hd__o2111ai_4 _24664_ (.A1(_14358_),
    .A2(_08006_),
    .B1(_05728_),
    .C1(_06154_),
    .D1(_08005_),
    .Y(_08009_));
 sky130_fd_sc_hd__nand2_4 _24665_ (.A(_08008_),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__xnor2_2 _24666_ (.A(_08004_),
    .B(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__xnor2_2 _24667_ (.A(_08003_),
    .B(_08011_),
    .Y(_08012_));
 sky130_vsdinv _24668_ (.A(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__nor2_1 _24669_ (.A(_07823_),
    .B(_07829_),
    .Y(_08014_));
 sky130_fd_sc_hd__o21bai_2 _24670_ (.A1(_07822_),
    .A2(_07830_),
    .B1_N(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__o21a_2 _24671_ (.A1(_06409_),
    .A2(_07825_),
    .B1(_07828_),
    .X(_08016_));
 sky130_fd_sc_hd__a2bb2oi_4 _24672_ (.A1_N(_14400_),
    .A2_N(_07850_),
    .B1(_07849_),
    .B2(_07851_),
    .Y(_08017_));
 sky130_fd_sc_hd__a22o_1 _24673_ (.A1(_06348_),
    .A2(_06040_),
    .B1(_06351_),
    .B2(_06412_),
    .X(_08018_));
 sky130_fd_sc_hd__nand3_4 _24674_ (.A(_06485_),
    .B(_06070_),
    .C(_05511_),
    .Y(_08019_));
 sky130_fd_sc_hd__or2b_1 _24675_ (.A(_08019_),
    .B_N(_05690_),
    .X(_08020_));
 sky130_fd_sc_hd__o2bb2ai_1 _24676_ (.A1_N(_08018_),
    .A2_N(_08020_),
    .B1(_14031_),
    .B2(_14372_),
    .Y(_08021_));
 sky130_fd_sc_hd__o2111ai_4 _24677_ (.A1(_06264_),
    .A2(_08019_),
    .B1(_06489_),
    .C1(_05699_),
    .D1(_08018_),
    .Y(_08022_));
 sky130_fd_sc_hd__nand2_4 _24678_ (.A(_08021_),
    .B(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__xnor2_4 _24679_ (.A(_08017_),
    .B(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__xor2_4 _24680_ (.A(_08016_),
    .B(_08024_),
    .X(_08025_));
 sky130_fd_sc_hd__xnor2_2 _24681_ (.A(_08015_),
    .B(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__nor2_4 _24682_ (.A(_08013_),
    .B(_08026_),
    .Y(_08027_));
 sky130_fd_sc_hd__nand2_1 _24683_ (.A(_08026_),
    .B(_08013_),
    .Y(_08028_));
 sky130_fd_sc_hd__nor3b_4 _24684_ (.A(_07998_),
    .B(_08027_),
    .C_N(_08028_),
    .Y(_08029_));
 sky130_vsdinv _24685_ (.A(_08029_),
    .Y(_08030_));
 sky130_vsdinv _24686_ (.A(_08027_),
    .Y(_08031_));
 sky130_fd_sc_hd__a21bo_1 _24687_ (.A1(_08031_),
    .A2(_08028_),
    .B1_N(_07998_),
    .X(_08032_));
 sky130_fd_sc_hd__nand2_1 _24688_ (.A(_08030_),
    .B(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__xor2_2 _24689_ (.A(_07997_),
    .B(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__nand2_2 _24690_ (.A(_07995_),
    .B(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__nand3b_4 _24691_ (.A_N(_08034_),
    .B(_07993_),
    .C(_07994_),
    .Y(_08036_));
 sky130_fd_sc_hd__nand3_4 _24692_ (.A(_07943_),
    .B(_08035_),
    .C(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__a21o_1 _24693_ (.A1(_08035_),
    .A2(_08036_),
    .B1(_07943_),
    .X(_08038_));
 sky130_vsdinv _24694_ (.A(_07768_),
    .Y(_08039_));
 sky130_fd_sc_hd__a21oi_4 _24695_ (.A1(_07767_),
    .A2(_07794_),
    .B1(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__nor2_1 _24696_ (.A(_07750_),
    .B(_07755_),
    .Y(_08041_));
 sky130_fd_sc_hd__o21ba_4 _24697_ (.A1(_07749_),
    .A2(_07756_),
    .B1_N(_08041_),
    .X(_08042_));
 sky130_fd_sc_hd__a2bb2oi_4 _24698_ (.A1_N(_14328_),
    .A2_N(_07752_),
    .B1(_07751_),
    .B2(_07753_),
    .Y(_08043_));
 sky130_fd_sc_hd__a2bb2oi_4 _24699_ (.A1_N(_14346_),
    .A2_N(_07805_),
    .B1(_07804_),
    .B2(_07806_),
    .Y(_08044_));
 sky130_fd_sc_hd__and2_2 _24700_ (.A(_04996_),
    .B(_06956_),
    .X(_08045_));
 sky130_fd_sc_hd__nand3_4 _24701_ (.A(_05486_),
    .B(_05063_),
    .C(\pcpi_mul.rs1[22] ),
    .Y(_08046_));
 sky130_fd_sc_hd__a22o_2 _24702_ (.A1(_05588_),
    .A2(\pcpi_mul.rs1[22] ),
    .B1(_05884_),
    .B2(\pcpi_mul.rs1[23] ),
    .X(_08047_));
 sky130_fd_sc_hd__o21ai_4 _24703_ (.A1(_14319_),
    .A2(_08046_),
    .B1(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__xor2_4 _24704_ (.A(_08045_),
    .B(_08048_),
    .X(_08049_));
 sky130_fd_sc_hd__xnor2_4 _24705_ (.A(_08044_),
    .B(_08049_),
    .Y(_08050_));
 sky130_fd_sc_hd__xor2_4 _24706_ (.A(_08043_),
    .B(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__nand3b_2 _24707_ (.A_N(_07816_),
    .B(_07813_),
    .C(_07812_),
    .Y(_08052_));
 sky130_fd_sc_hd__or2b_1 _24708_ (.A(_07817_),
    .B_N(_07808_),
    .X(_08053_));
 sky130_fd_sc_hd__nand3b_2 _24709_ (.A_N(_08051_),
    .B(_08052_),
    .C(_08053_),
    .Y(_08054_));
 sky130_fd_sc_hd__nand2_1 _24710_ (.A(_08053_),
    .B(_08052_),
    .Y(_08055_));
 sky130_fd_sc_hd__nand2_2 _24711_ (.A(_08055_),
    .B(_08051_),
    .Y(_08056_));
 sky130_fd_sc_hd__nand2_4 _24712_ (.A(_08054_),
    .B(_08056_),
    .Y(_08057_));
 sky130_fd_sc_hd__nor2_1 _24713_ (.A(_08042_),
    .B(_08057_),
    .Y(_08058_));
 sky130_vsdinv _24714_ (.A(_08058_),
    .Y(_08059_));
 sky130_fd_sc_hd__nand2_2 _24715_ (.A(_08057_),
    .B(_08042_),
    .Y(_08060_));
 sky130_fd_sc_hd__and2_1 _24716_ (.A(_07759_),
    .B(_07757_),
    .X(_08061_));
 sky130_fd_sc_hd__a211o_2 _24717_ (.A1(_08059_),
    .A2(_08060_),
    .B1(_08061_),
    .C1(_07764_),
    .X(_08062_));
 sky130_fd_sc_hd__o211ai_4 _24718_ (.A1(_08061_),
    .A2(_07764_),
    .B1(_08059_),
    .C1(_08060_),
    .Y(_08063_));
 sky130_fd_sc_hd__clkbuf_4 _24719_ (.A(_07585_),
    .X(_08064_));
 sky130_fd_sc_hd__buf_4 _24720_ (.A(_08064_),
    .X(_08065_));
 sky130_fd_sc_hd__nor3_4 _24721_ (.A(_06433_),
    .B(_14305_),
    .C(_07780_),
    .Y(_08066_));
 sky130_fd_sc_hd__a41oi_4 _24722_ (.A1(_05403_),
    .A2(_05899_),
    .A3(_08065_),
    .A4(_07770_),
    .B1(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__nor2_1 _24723_ (.A(_07783_),
    .B(_07790_),
    .Y(_08068_));
 sky130_fd_sc_hd__o21bai_4 _24724_ (.A1(_07781_),
    .A2(_07791_),
    .B1_N(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__buf_2 _24725_ (.A(_07485_),
    .X(_08070_));
 sky130_fd_sc_hd__and2_2 _24726_ (.A(_06025_),
    .B(_08070_),
    .X(_08071_));
 sky130_fd_sc_hd__nand2_2 _24727_ (.A(_04936_),
    .B(_07585_),
    .Y(_08072_));
 sky130_fd_sc_hd__clkbuf_4 _24728_ (.A(\pcpi_mul.rs1[29] ),
    .X(_08073_));
 sky130_fd_sc_hd__nand2_2 _24729_ (.A(_04938_),
    .B(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__xnor2_4 _24730_ (.A(_08072_),
    .B(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__xor2_4 _24731_ (.A(_08071_),
    .B(_08075_),
    .X(_08076_));
 sky130_fd_sc_hd__buf_2 _24732_ (.A(\pcpi_mul.rs1[30] ),
    .X(_08077_));
 sky130_fd_sc_hd__buf_2 _24733_ (.A(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__and2_2 _24734_ (.A(_04955_),
    .B(_08078_),
    .X(_08079_));
 sky130_fd_sc_hd__nand3_4 _24735_ (.A(_05419_),
    .B(_05324_),
    .C(_07044_),
    .Y(_08080_));
 sky130_fd_sc_hd__a22o_2 _24736_ (.A1(_05116_),
    .A2(_07209_),
    .B1(_06445_),
    .B2(_07476_),
    .X(_08081_));
 sky130_fd_sc_hd__o21ai_4 _24737_ (.A1(_14303_),
    .A2(_08080_),
    .B1(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__xor2_4 _24738_ (.A(_08079_),
    .B(_08082_),
    .X(_08083_));
 sky130_fd_sc_hd__buf_4 _24739_ (.A(_14285_),
    .X(_08084_));
 sky130_fd_sc_hd__buf_2 _24740_ (.A(_06957_),
    .X(_08085_));
 sky130_fd_sc_hd__nand3b_1 _24741_ (.A_N(_07787_),
    .B(_06159_),
    .C(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__o31a_2 _24742_ (.A1(_14097_),
    .A2(_08084_),
    .A3(_07789_),
    .B1(_08086_),
    .X(_08087_));
 sky130_fd_sc_hd__xnor2_4 _24743_ (.A(_08083_),
    .B(_08087_),
    .Y(_08088_));
 sky130_fd_sc_hd__xor2_4 _24744_ (.A(_08076_),
    .B(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__xnor2_4 _24745_ (.A(_08069_),
    .B(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__xor2_4 _24746_ (.A(_08067_),
    .B(_08090_),
    .X(_08091_));
 sky130_fd_sc_hd__a21o_2 _24747_ (.A1(_08062_),
    .A2(_08063_),
    .B1(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__nand3_4 _24748_ (.A(_08062_),
    .B(_08091_),
    .C(_08063_),
    .Y(_08093_));
 sky130_fd_sc_hd__a21o_2 _24749_ (.A1(_07843_),
    .A2(_07841_),
    .B1(_07838_),
    .X(_08094_));
 sky130_fd_sc_hd__a21oi_4 _24750_ (.A1(_08092_),
    .A2(_08093_),
    .B1(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__nand3_4 _24751_ (.A(_08092_),
    .B(_08094_),
    .C(_08093_),
    .Y(_08096_));
 sky130_fd_sc_hd__nor3b_4 _24752_ (.A(_08040_),
    .B(_08095_),
    .C_N(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__and3_1 _24753_ (.A(_08092_),
    .B(_08094_),
    .C(_08093_),
    .X(_08098_));
 sky130_fd_sc_hd__o21a_1 _24754_ (.A1(_08095_),
    .A2(_08098_),
    .B1(_08040_),
    .X(_08099_));
 sky130_fd_sc_hd__o2bb2ai_2 _24755_ (.A1_N(_08037_),
    .A2_N(_08038_),
    .B1(_08097_),
    .B2(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__nor2_2 _24756_ (.A(_08097_),
    .B(_08099_),
    .Y(_08101_));
 sky130_fd_sc_hd__nand3_4 _24757_ (.A(_08038_),
    .B(_08101_),
    .C(_08037_),
    .Y(_08102_));
 sky130_fd_sc_hd__nand2_1 _24758_ (.A(_08100_),
    .B(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__o21ba_1 _24759_ (.A1(_07899_),
    .A2(_07901_),
    .B1_N(_07902_),
    .X(_08104_));
 sky130_fd_sc_hd__o21a_1 _24760_ (.A1(_07907_),
    .A2(_08104_),
    .B1(_07905_),
    .X(_08105_));
 sky130_fd_sc_hd__nand2_2 _24761_ (.A(_08103_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__o21ai_2 _24762_ (.A1(_07907_),
    .A2(_08104_),
    .B1(_07905_),
    .Y(_08107_));
 sky130_fd_sc_hd__nand3_4 _24763_ (.A(_08107_),
    .B(_08102_),
    .C(_08100_),
    .Y(_08108_));
 sky130_fd_sc_hd__nor2_1 _24764_ (.A(_07772_),
    .B(_07793_),
    .Y(_08109_));
 sky130_fd_sc_hd__a21o_4 _24765_ (.A1(_07792_),
    .A2(_07774_),
    .B1(_08109_),
    .X(_08110_));
 sky130_fd_sc_hd__a21boi_4 _24766_ (.A1(_07798_),
    .A2(_07801_),
    .B1_N(_07799_),
    .Y(_08111_));
 sky130_fd_sc_hd__xnor2_4 _24767_ (.A(_08110_),
    .B(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__a21oi_2 _24768_ (.A1(_08106_),
    .A2(_08108_),
    .B1(_08112_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand3_4 _24769_ (.A(_08106_),
    .B(_08112_),
    .C(_08108_),
    .Y(_08114_));
 sky130_vsdinv _24770_ (.A(_08114_),
    .Y(_08115_));
 sky130_vsdinv _24771_ (.A(_07920_),
    .Y(_08116_));
 sky130_fd_sc_hd__a21oi_2 _24772_ (.A1(_07913_),
    .A2(_07914_),
    .B1(_07912_),
    .Y(_08117_));
 sky130_fd_sc_hd__o21ai_4 _24773_ (.A1(_08116_),
    .A2(_08117_),
    .B1(_07915_),
    .Y(_08118_));
 sky130_fd_sc_hd__o21bai_4 _24774_ (.A1(_08113_),
    .A2(_08115_),
    .B1_N(_08118_),
    .Y(_08119_));
 sky130_fd_sc_hd__a21o_1 _24775_ (.A1(_08106_),
    .A2(_08108_),
    .B1(_08112_),
    .X(_08120_));
 sky130_fd_sc_hd__nand3_4 _24776_ (.A(_08120_),
    .B(_08118_),
    .C(_08114_),
    .Y(_08121_));
 sky130_fd_sc_hd__a21oi_1 _24777_ (.A1(_08119_),
    .A2(_08121_),
    .B1(_07928_),
    .Y(_08122_));
 sky130_fd_sc_hd__nand3_4 _24778_ (.A(_08119_),
    .B(_07928_),
    .C(_08121_),
    .Y(_08123_));
 sky130_vsdinv _24779_ (.A(_08123_),
    .Y(_08124_));
 sky130_vsdinv _24780_ (.A(_07712_),
    .Y(_08125_));
 sky130_fd_sc_hd__o21ai_4 _24781_ (.A1(_08125_),
    .A2(_07936_),
    .B1(_07930_),
    .Y(_08126_));
 sky130_fd_sc_hd__o21bai_2 _24782_ (.A1(_08122_),
    .A2(_08124_),
    .B1_N(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__a21o_1 _24783_ (.A1(_08119_),
    .A2(_08121_),
    .B1(_07928_),
    .X(_08128_));
 sky130_fd_sc_hd__nand3_4 _24784_ (.A(_08128_),
    .B(_08123_),
    .C(_08126_),
    .Y(_08129_));
 sky130_fd_sc_hd__nand2_4 _24785_ (.A(_08127_),
    .B(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__nand2_1 _24786_ (.A(_07730_),
    .B(_07733_),
    .Y(_08131_));
 sky130_fd_sc_hd__nor2_4 _24787_ (.A(_08131_),
    .B(_07940_),
    .Y(_08132_));
 sky130_fd_sc_hd__a21oi_4 _24788_ (.A1(_07938_),
    .A2(_07932_),
    .B1(_07934_),
    .Y(_08133_));
 sky130_fd_sc_hd__a21oi_4 _24789_ (.A1(_07733_),
    .A2(_07939_),
    .B1(_08133_),
    .Y(_08134_));
 sky130_fd_sc_hd__a21oi_4 _24790_ (.A1(_07745_),
    .A2(_08132_),
    .B1(_08134_),
    .Y(_08135_));
 sky130_fd_sc_hd__xor2_4 _24791_ (.A(_08130_),
    .B(_08135_),
    .X(_02649_));
 sky130_fd_sc_hd__nor2_1 _24792_ (.A(_08044_),
    .B(_08049_),
    .Y(_08136_));
 sky130_fd_sc_hd__o21ba_2 _24793_ (.A1(_08043_),
    .A2(_08050_),
    .B1_N(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__or2b_1 _24794_ (.A(_08011_),
    .B_N(_08003_),
    .X(_08138_));
 sky130_fd_sc_hd__o21ai_2 _24795_ (.A1(_08010_),
    .A2(_08004_),
    .B1(_08138_),
    .Y(_08139_));
 sky130_fd_sc_hd__a2bb2oi_4 _24796_ (.A1_N(_14321_),
    .A2_N(_08046_),
    .B1(_08045_),
    .B2(_08047_),
    .Y(_08140_));
 sky130_fd_sc_hd__a2bb2oi_4 _24797_ (.A1_N(_14339_),
    .A2_N(_08000_),
    .B1(_07999_),
    .B2(_08001_),
    .Y(_08141_));
 sky130_fd_sc_hd__and2_2 _24798_ (.A(_06001_),
    .B(_07786_),
    .X(_08142_));
 sky130_fd_sc_hd__nand3_4 _24799_ (.A(_14062_),
    .B(_05163_),
    .C(_07204_),
    .Y(_08143_));
 sky130_fd_sc_hd__a22o_2 _24800_ (.A1(_05486_),
    .A2(\pcpi_mul.rs1[23] ),
    .B1(_14066_),
    .B2(\pcpi_mul.rs1[24] ),
    .X(_08144_));
 sky130_fd_sc_hd__o21ai_4 _24801_ (.A1(_14313_),
    .A2(_08143_),
    .B1(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__xor2_4 _24802_ (.A(_08142_),
    .B(_08145_),
    .X(_08146_));
 sky130_fd_sc_hd__xnor2_4 _24803_ (.A(_08141_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__xor2_4 _24804_ (.A(_08140_),
    .B(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__xnor2_1 _24805_ (.A(_08139_),
    .B(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__nor2_2 _24806_ (.A(_08137_),
    .B(_08149_),
    .Y(_08150_));
 sky130_vsdinv _24807_ (.A(_08150_),
    .Y(_08151_));
 sky130_fd_sc_hd__nand2_2 _24808_ (.A(_08149_),
    .B(_08137_),
    .Y(_08152_));
 sky130_fd_sc_hd__o21ai_4 _24809_ (.A1(_08042_),
    .A2(_08057_),
    .B1(_08056_),
    .Y(_08153_));
 sky130_fd_sc_hd__a21o_2 _24810_ (.A1(_08151_),
    .A2(_08152_),
    .B1(_08153_),
    .X(_08154_));
 sky130_fd_sc_hd__nand3b_4 _24811_ (.A_N(_08150_),
    .B(_08152_),
    .C(_08153_),
    .Y(_08155_));
 sky130_fd_sc_hd__nand2_1 _24812_ (.A(_08154_),
    .B(_08155_),
    .Y(_08156_));
 sky130_fd_sc_hd__clkbuf_2 _24813_ (.A(_08073_),
    .X(_08157_));
 sky130_fd_sc_hd__buf_4 _24814_ (.A(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__nor3_4 _24815_ (.A(_06433_),
    .B(_14300_),
    .C(_08075_),
    .Y(_08159_));
 sky130_fd_sc_hd__a41oi_4 _24816_ (.A1(_05298_),
    .A2(_05899_),
    .A3(_08158_),
    .A4(_08065_),
    .B1(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__nor2_1 _24817_ (.A(_08083_),
    .B(_08087_),
    .Y(_08161_));
 sky130_fd_sc_hd__o21bai_4 _24818_ (.A1(_08076_),
    .A2(_08088_),
    .B1_N(_08161_),
    .Y(_08162_));
 sky130_fd_sc_hd__and2_2 _24819_ (.A(_06025_),
    .B(_07778_),
    .X(_08163_));
 sky130_fd_sc_hd__nand2_2 _24820_ (.A(_04884_),
    .B(_08073_),
    .Y(_08164_));
 sky130_fd_sc_hd__buf_2 _24821_ (.A(_08077_),
    .X(_08165_));
 sky130_fd_sc_hd__nand2_2 _24822_ (.A(_04876_),
    .B(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__xnor2_4 _24823_ (.A(_08164_),
    .B(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__xor2_4 _24824_ (.A(_08163_),
    .B(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__a2bb2oi_4 _24825_ (.A1_N(_14304_),
    .A2_N(_08080_),
    .B1(_08079_),
    .B2(_08081_),
    .Y(_08169_));
 sky130_fd_sc_hd__clkbuf_2 _24826_ (.A(\pcpi_mul.rs1[31] ),
    .X(_08170_));
 sky130_fd_sc_hd__buf_2 _24827_ (.A(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__nand2_4 _24828_ (.A(_05319_),
    .B(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__or4_4 _24829_ (.A(_14074_),
    .B(_14077_),
    .C(_14296_),
    .D(_14302_),
    .X(_08173_));
 sky130_fd_sc_hd__a22o_1 _24830_ (.A1(_05116_),
    .A2(_07476_),
    .B1(_06445_),
    .B2(_07484_),
    .X(_08174_));
 sky130_fd_sc_hd__nand2_2 _24831_ (.A(_08173_),
    .B(_08174_),
    .Y(_08175_));
 sky130_fd_sc_hd__xnor2_4 _24832_ (.A(_08172_),
    .B(_08175_),
    .Y(_08176_));
 sky130_fd_sc_hd__xnor2_4 _24833_ (.A(_08169_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__xor2_4 _24834_ (.A(_08168_),
    .B(_08177_),
    .X(_08178_));
 sky130_fd_sc_hd__xnor2_4 _24835_ (.A(_08162_),
    .B(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__xor2_4 _24836_ (.A(_08160_),
    .B(_08179_),
    .X(_08180_));
 sky130_fd_sc_hd__and2b_1 _24837_ (.A_N(_08156_),
    .B(_08180_),
    .X(_08181_));
 sky130_vsdinv _24838_ (.A(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__a21o_1 _24839_ (.A1(_08155_),
    .A2(_08154_),
    .B1(_08180_),
    .X(_08183_));
 sky130_fd_sc_hd__a21o_1 _24840_ (.A1(_08032_),
    .A2(_07997_),
    .B1(_08029_),
    .X(_08184_));
 sky130_fd_sc_hd__a21o_1 _24841_ (.A1(_08182_),
    .A2(_08183_),
    .B1(_08184_),
    .X(_08185_));
 sky130_fd_sc_hd__nand3b_4 _24842_ (.A_N(_08181_),
    .B(_08184_),
    .C(_08183_),
    .Y(_08186_));
 sky130_fd_sc_hd__a21boi_1 _24843_ (.A1(_08062_),
    .A2(_08091_),
    .B1_N(_08063_),
    .Y(_08187_));
 sky130_vsdinv _24844_ (.A(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__a21oi_4 _24845_ (.A1(_08185_),
    .A2(_08186_),
    .B1(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__nand3_4 _24846_ (.A(_08185_),
    .B(_08188_),
    .C(_08186_),
    .Y(_08190_));
 sky130_vsdinv _24847_ (.A(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__nor2_4 _24848_ (.A(_08189_),
    .B(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__and2_2 _24849_ (.A(_05720_),
    .B(_07033_),
    .X(_08193_));
 sky130_fd_sc_hd__nand3_4 _24850_ (.A(_05582_),
    .B(_05273_),
    .C(_06577_),
    .Y(_08194_));
 sky130_fd_sc_hd__a22o_2 _24851_ (.A1(_05359_),
    .A2(_07746_),
    .B1(_05363_),
    .B2(_06587_),
    .X(_08195_));
 sky130_fd_sc_hd__o21ai_4 _24852_ (.A1(_07214_),
    .A2(_08194_),
    .B1(_08195_),
    .Y(_08196_));
 sky130_fd_sc_hd__xnor2_4 _24853_ (.A(_08193_),
    .B(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__o21a_4 _24854_ (.A1(_14359_),
    .A2(_08006_),
    .B1(_08009_),
    .X(_08198_));
 sky130_fd_sc_hd__clkbuf_4 _24855_ (.A(_05732_),
    .X(_08199_));
 sky130_fd_sc_hd__a22o_1 _24856_ (.A1(_05955_),
    .A2(_06028_),
    .B1(_08199_),
    .B2(_06287_),
    .X(_08200_));
 sky130_fd_sc_hd__nand3_4 _24857_ (.A(_14036_),
    .B(_14041_),
    .C(_06028_),
    .Y(_08201_));
 sky130_fd_sc_hd__or2b_1 _24858_ (.A(_08201_),
    .B_N(_06154_),
    .X(_08202_));
 sky130_fd_sc_hd__o2bb2ai_2 _24859_ (.A1_N(_08200_),
    .A2_N(_08202_),
    .B1(_06207_),
    .B2(_14346_),
    .Y(_08203_));
 sky130_fd_sc_hd__o2111ai_4 _24860_ (.A1(_14352_),
    .A2(_08201_),
    .B1(_05441_),
    .C1(_06165_),
    .D1(_08200_),
    .Y(_08204_));
 sky130_fd_sc_hd__nand2_4 _24861_ (.A(_08203_),
    .B(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__xnor2_4 _24862_ (.A(_08198_),
    .B(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__xor2_4 _24863_ (.A(_08197_),
    .B(_08206_),
    .X(_08207_));
 sky130_fd_sc_hd__nor2_1 _24864_ (.A(_08017_),
    .B(_08023_),
    .Y(_08208_));
 sky130_fd_sc_hd__o21bai_2 _24865_ (.A1(_08016_),
    .A2(_08024_),
    .B1_N(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__buf_6 _24866_ (.A(_14378_),
    .X(_08210_));
 sky130_fd_sc_hd__o21a_4 _24867_ (.A1(_08210_),
    .A2(_08019_),
    .B1(_08022_),
    .X(_08211_));
 sky130_fd_sc_hd__a2bb2oi_4 _24868_ (.A1_N(_14394_),
    .A2_N(_07974_),
    .B1(_07973_),
    .B2(_07975_),
    .Y(_08212_));
 sky130_fd_sc_hd__a22o_1 _24869_ (.A1(_14023_),
    .A2(_06412_),
    .B1(_14027_),
    .B2(_05698_),
    .X(_08213_));
 sky130_fd_sc_hd__nand3_4 _24870_ (.A(_06348_),
    .B(_06070_),
    .C(_14376_),
    .Y(_08214_));
 sky130_fd_sc_hd__or2b_1 _24871_ (.A(_08214_),
    .B_N(_05768_),
    .X(_08215_));
 sky130_fd_sc_hd__o2bb2ai_1 _24872_ (.A1_N(_08213_),
    .A2_N(_08215_),
    .B1(_14031_),
    .B2(_14366_),
    .Y(_08216_));
 sky130_fd_sc_hd__o2111ai_4 _24873_ (.A1(_14371_),
    .A2(_08214_),
    .B1(_06355_),
    .C1(_05777_),
    .D1(_08213_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2_4 _24874_ (.A(_08216_),
    .B(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__xnor2_4 _24875_ (.A(_08212_),
    .B(_08218_),
    .Y(_08219_));
 sky130_fd_sc_hd__xor2_4 _24876_ (.A(_08211_),
    .B(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__xnor2_2 _24877_ (.A(_08209_),
    .B(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__nor2_2 _24878_ (.A(_08207_),
    .B(_08221_),
    .Y(_08222_));
 sky130_fd_sc_hd__and2_1 _24879_ (.A(_08221_),
    .B(_08207_),
    .X(_08223_));
 sky130_fd_sc_hd__and2_1 _24880_ (.A(_07987_),
    .B(_07972_),
    .X(_08224_));
 sky130_fd_sc_hd__o21bai_1 _24881_ (.A1(_07970_),
    .A2(_07988_),
    .B1_N(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__or3b_4 _24882_ (.A(_08222_),
    .B(_08223_),
    .C_N(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__o21bai_2 _24883_ (.A1(_08222_),
    .A2(_08223_),
    .B1_N(_08225_),
    .Y(_08227_));
 sky130_fd_sc_hd__a21oi_1 _24884_ (.A1(_08025_),
    .A2(_08015_),
    .B1(_08027_),
    .Y(_08228_));
 sky130_fd_sc_hd__a21bo_1 _24885_ (.A1(_08226_),
    .A2(_08227_),
    .B1_N(_08228_),
    .X(_08229_));
 sky130_fd_sc_hd__nand3b_4 _24886_ (.A_N(_08228_),
    .B(_08226_),
    .C(_08227_),
    .Y(_08230_));
 sky130_fd_sc_hd__nand2_2 _24887_ (.A(_08229_),
    .B(_08230_),
    .Y(_08231_));
 sky130_vsdinv _24888_ (.A(_07968_),
    .Y(_08232_));
 sky130_fd_sc_hd__a21oi_2 _24889_ (.A1(_08232_),
    .A2(_07989_),
    .B1(_07967_),
    .Y(_08233_));
 sky130_fd_sc_hd__nand2_1 _24890_ (.A(_07959_),
    .B(_07957_),
    .Y(_08234_));
 sky130_fd_sc_hd__o21a_2 _24891_ (.A1(_07948_),
    .A2(_07951_),
    .B1(_07949_),
    .X(_08235_));
 sky130_fd_sc_hd__a22o_1 _24892_ (.A1(_07264_),
    .A2(_04978_),
    .B1(_07265_),
    .B2(_05091_),
    .X(_08236_));
 sky130_fd_sc_hd__nand3_4 _24893_ (.A(_07264_),
    .B(_07265_),
    .C(_05959_),
    .Y(_08237_));
 sky130_fd_sc_hd__or2b_1 _24894_ (.A(_08237_),
    .B_N(_05099_),
    .X(_08238_));
 sky130_fd_sc_hd__o2bb2ai_1 _24895_ (.A1_N(_08236_),
    .A2_N(_08238_),
    .B1(_13993_),
    .B2(_05115_),
    .Y(_08239_));
 sky130_fd_sc_hd__o2111ai_4 _24896_ (.A1(_05057_),
    .A2(_08237_),
    .B1(_07106_),
    .C1(_05819_),
    .D1(_08236_),
    .Y(_08240_));
 sky130_fd_sc_hd__nand2_2 _24897_ (.A(_08239_),
    .B(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__xnor2_2 _24898_ (.A(_08235_),
    .B(_08241_),
    .Y(_08242_));
 sky130_fd_sc_hd__xor2_2 _24899_ (.A(_08234_),
    .B(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__buf_6 _24900_ (.A(_07946_),
    .X(_08244_));
 sky130_fd_sc_hd__nand3b_4 _24901_ (.A_N(_07952_),
    .B(_08244_),
    .C(_04719_),
    .Y(_08245_));
 sky130_fd_sc_hd__nand2_2 _24902_ (.A(_13961_),
    .B(_05533_),
    .Y(_08246_));
 sky130_fd_sc_hd__nand2_2 _24903_ (.A(_07945_),
    .B(_04872_),
    .Y(_08247_));
 sky130_fd_sc_hd__xnor2_4 _24904_ (.A(_08246_),
    .B(_08247_),
    .Y(_08248_));
 sky130_fd_sc_hd__and2_2 _24905_ (.A(\pcpi_mul.rs2[27] ),
    .B(_04976_),
    .X(_08249_));
 sky130_fd_sc_hd__nand2_2 _24906_ (.A(_13976_),
    .B(_04949_),
    .Y(_08250_));
 sky130_fd_sc_hd__and2_1 _24907_ (.A(\pcpi_mul.rs2[29] ),
    .B(_04889_),
    .X(_08251_));
 sky130_fd_sc_hd__xor2_4 _24908_ (.A(_08250_),
    .B(_08251_),
    .X(_08252_));
 sky130_fd_sc_hd__xor2_4 _24909_ (.A(_08249_),
    .B(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__xnor2_2 _24910_ (.A(_08248_),
    .B(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__xor2_2 _24911_ (.A(_08245_),
    .B(_08254_),
    .X(_08255_));
 sky130_fd_sc_hd__xor2_1 _24912_ (.A(_08243_),
    .B(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__a21bo_1 _24913_ (.A1(_07953_),
    .A2(_07965_),
    .B1_N(_08256_),
    .X(_08257_));
 sky130_fd_sc_hd__nand3b_2 _24914_ (.A_N(_08256_),
    .B(_07953_),
    .C(_07965_),
    .Y(_08258_));
 sky130_fd_sc_hd__nor2_1 _24915_ (.A(_07978_),
    .B(_07985_),
    .Y(_08259_));
 sky130_fd_sc_hd__o21ba_1 _24916_ (.A1(_07977_),
    .A2(_07986_),
    .B1_N(_08259_),
    .X(_08260_));
 sky130_fd_sc_hd__buf_2 _24917_ (.A(_06319_),
    .X(_08261_));
 sky130_fd_sc_hd__and2_2 _24918_ (.A(_08261_),
    .B(_06160_),
    .X(_08262_));
 sky130_fd_sc_hd__nand3_4 _24919_ (.A(_06895_),
    .B(_14015_),
    .C(_05322_),
    .Y(_08263_));
 sky130_fd_sc_hd__buf_2 _24920_ (.A(_05917_),
    .X(_08264_));
 sky130_fd_sc_hd__a22o_2 _24921_ (.A1(_14010_),
    .A2(_05497_),
    .B1(_06185_),
    .B2(_08264_),
    .X(_08265_));
 sky130_fd_sc_hd__o21ai_4 _24922_ (.A1(_14389_),
    .A2(_08263_),
    .B1(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__xor2_4 _24923_ (.A(_08262_),
    .B(_08266_),
    .X(_08267_));
 sky130_fd_sc_hd__o21a_2 _24924_ (.A1(_14411_),
    .A2(_07981_),
    .B1(_07984_),
    .X(_08268_));
 sky130_fd_sc_hd__buf_4 _24925_ (.A(_13997_),
    .X(_08269_));
 sky130_fd_sc_hd__a22o_1 _24926_ (.A1(_08269_),
    .A2(_05427_),
    .B1(_07979_),
    .B2(_05181_),
    .X(_08270_));
 sky130_fd_sc_hd__nand3_4 _24927_ (.A(_06744_),
    .B(_14001_),
    .C(_05227_),
    .Y(_08271_));
 sky130_fd_sc_hd__or2b_1 _24928_ (.A(_08271_),
    .B_N(_05516_),
    .X(_08272_));
 sky130_fd_sc_hd__o2bb2ai_1 _24929_ (.A1_N(_08270_),
    .A2_N(_08272_),
    .B1(_14005_),
    .B2(_14400_),
    .Y(_08273_));
 sky130_fd_sc_hd__o2111ai_4 _24930_ (.A1(_06127_),
    .A2(_08271_),
    .B1(_06470_),
    .C1(_05405_),
    .D1(_08270_),
    .Y(_08274_));
 sky130_fd_sc_hd__nand2_4 _24931_ (.A(_08273_),
    .B(_08274_),
    .Y(_08275_));
 sky130_fd_sc_hd__xnor2_4 _24932_ (.A(_08268_),
    .B(_08275_),
    .Y(_08276_));
 sky130_fd_sc_hd__xor2_4 _24933_ (.A(_08267_),
    .B(_08276_),
    .X(_08277_));
 sky130_fd_sc_hd__a21o_1 _24934_ (.A1(_07883_),
    .A2(_07885_),
    .B1(_07964_),
    .X(_08278_));
 sky130_fd_sc_hd__o21ai_2 _24935_ (.A1(_07963_),
    .A2(_07960_),
    .B1(_08278_),
    .Y(_08279_));
 sky130_fd_sc_hd__xnor2_2 _24936_ (.A(_08277_),
    .B(_08279_),
    .Y(_08280_));
 sky130_fd_sc_hd__xor2_2 _24937_ (.A(_08260_),
    .B(_08280_),
    .X(_08281_));
 sky130_fd_sc_hd__a21oi_2 _24938_ (.A1(_08257_),
    .A2(_08258_),
    .B1(_08281_),
    .Y(_08282_));
 sky130_fd_sc_hd__and3_1 _24939_ (.A(_08257_),
    .B(_08281_),
    .C(_08258_),
    .X(_08283_));
 sky130_fd_sc_hd__or3_4 _24940_ (.A(_08233_),
    .B(_08282_),
    .C(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__o21ai_2 _24941_ (.A1(_08282_),
    .A2(_08283_),
    .B1(_08233_),
    .Y(_08285_));
 sky130_fd_sc_hd__nand2_2 _24942_ (.A(_08284_),
    .B(_08285_),
    .Y(_08286_));
 sky130_fd_sc_hd__nor2_4 _24943_ (.A(_08231_),
    .B(_08286_),
    .Y(_08287_));
 sky130_fd_sc_hd__nand2_1 _24944_ (.A(_08036_),
    .B(_07993_),
    .Y(_08288_));
 sky130_fd_sc_hd__a22oi_4 _24945_ (.A1(_08230_),
    .A2(_08229_),
    .B1(_08284_),
    .B2(_08285_),
    .Y(_08289_));
 sky130_vsdinv _24946_ (.A(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__nand3b_4 _24947_ (.A_N(_08287_),
    .B(_08288_),
    .C(_08290_),
    .Y(_08291_));
 sky130_fd_sc_hd__o211ai_4 _24948_ (.A1(_08289_),
    .A2(_08287_),
    .B1(_07993_),
    .C1(_08036_),
    .Y(_08292_));
 sky130_fd_sc_hd__nand3_4 _24949_ (.A(_08192_),
    .B(_08291_),
    .C(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__o2bb2ai_2 _24950_ (.A1_N(_08291_),
    .A2_N(_08292_),
    .B1(_08191_),
    .B2(_08189_),
    .Y(_08294_));
 sky130_fd_sc_hd__nand2_2 _24951_ (.A(_08102_),
    .B(_08037_),
    .Y(_08295_));
 sky130_fd_sc_hd__a21oi_1 _24952_ (.A1(_08293_),
    .A2(_08294_),
    .B1(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__nand3_4 _24953_ (.A(_08295_),
    .B(_08293_),
    .C(_08294_),
    .Y(_08297_));
 sky130_vsdinv _24954_ (.A(_08297_),
    .Y(_08298_));
 sky130_fd_sc_hd__nor2_1 _24955_ (.A(_08067_),
    .B(_08090_),
    .Y(_08299_));
 sky130_fd_sc_hd__a21o_4 _24956_ (.A1(_08089_),
    .A2(_08069_),
    .B1(_08299_),
    .X(_08300_));
 sky130_fd_sc_hd__o21ai_4 _24957_ (.A1(_08040_),
    .A2(_08095_),
    .B1(_08096_),
    .Y(_08301_));
 sky130_fd_sc_hd__xor2_4 _24958_ (.A(_08300_),
    .B(_08301_),
    .X(_08302_));
 sky130_fd_sc_hd__o21bai_2 _24959_ (.A1(_08296_),
    .A2(_08298_),
    .B1_N(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__a21o_1 _24960_ (.A1(_08293_),
    .A2(_08294_),
    .B1(_08295_),
    .X(_08304_));
 sky130_fd_sc_hd__nand3_4 _24961_ (.A(_08304_),
    .B(_08302_),
    .C(_08297_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_1 _24962_ (.A(_08303_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__nand2_2 _24963_ (.A(_08114_),
    .B(_08108_),
    .Y(_08307_));
 sky130_vsdinv _24964_ (.A(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__nand2_2 _24965_ (.A(_08306_),
    .B(_08308_),
    .Y(_08309_));
 sky130_fd_sc_hd__nand3_4 _24966_ (.A(_08303_),
    .B(_08307_),
    .C(_08305_),
    .Y(_08310_));
 sky130_fd_sc_hd__a21boi_4 _24967_ (.A1(_07803_),
    .A2(_07799_),
    .B1_N(_08110_),
    .Y(_08311_));
 sky130_fd_sc_hd__a21o_1 _24968_ (.A1(_08309_),
    .A2(_08310_),
    .B1(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__nand3_4 _24969_ (.A(_08309_),
    .B(_08311_),
    .C(_08310_),
    .Y(_08313_));
 sky130_vsdinv _24970_ (.A(_07928_),
    .Y(_08314_));
 sky130_fd_sc_hd__a21oi_2 _24971_ (.A1(_08120_),
    .A2(_08114_),
    .B1(_08118_),
    .Y(_08315_));
 sky130_fd_sc_hd__o21ai_4 _24972_ (.A1(_08314_),
    .A2(_08315_),
    .B1(_08121_),
    .Y(_08316_));
 sky130_fd_sc_hd__a21oi_4 _24973_ (.A1(_08312_),
    .A2(_08313_),
    .B1(_08316_),
    .Y(_08317_));
 sky130_fd_sc_hd__a21boi_2 _24974_ (.A1(_08119_),
    .A2(_07928_),
    .B1_N(_08121_),
    .Y(_08318_));
 sky130_fd_sc_hd__a21oi_4 _24975_ (.A1(_08309_),
    .A2(_08310_),
    .B1(_08311_),
    .Y(_08319_));
 sky130_vsdinv _24976_ (.A(_08313_),
    .Y(_08320_));
 sky130_fd_sc_hd__nor3_4 _24977_ (.A(_08318_),
    .B(_08319_),
    .C(_08320_),
    .Y(_08321_));
 sky130_fd_sc_hd__nor2_8 _24978_ (.A(_08317_),
    .B(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__a21oi_4 _24979_ (.A1(_08128_),
    .A2(_08123_),
    .B1(_08126_),
    .Y(_08323_));
 sky130_vsdinv _24980_ (.A(_08129_),
    .Y(_08324_));
 sky130_fd_sc_hd__o21bai_4 _24981_ (.A1(_08323_),
    .A2(_08135_),
    .B1_N(_08324_),
    .Y(_08325_));
 sky130_fd_sc_hd__xor2_4 _24982_ (.A(_08322_),
    .B(_08325_),
    .X(_02650_));
 sky130_fd_sc_hd__and2_1 _24983_ (.A(_08220_),
    .B(_08209_),
    .X(_08326_));
 sky130_fd_sc_hd__o21ba_1 _24984_ (.A1(_08207_),
    .A2(_08221_),
    .B1_N(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__nand2_1 _24985_ (.A(_08279_),
    .B(_08277_),
    .Y(_08328_));
 sky130_fd_sc_hd__o21a_1 _24986_ (.A1(_08260_),
    .A2(_08280_),
    .B1(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__clkbuf_4 _24987_ (.A(_07027_),
    .X(_08330_));
 sky130_fd_sc_hd__and2_2 _24988_ (.A(_05206_),
    .B(_08330_),
    .X(_08331_));
 sky130_fd_sc_hd__buf_6 _24989_ (.A(_14327_),
    .X(_08332_));
 sky130_fd_sc_hd__buf_4 _24990_ (.A(_05359_),
    .X(_08333_));
 sky130_fd_sc_hd__nand3_4 _24991_ (.A(_08333_),
    .B(_05274_),
    .C(_07481_),
    .Y(_08334_));
 sky130_fd_sc_hd__a22o_2 _24992_ (.A1(_08333_),
    .A2(_07481_),
    .B1(_05274_),
    .B2(_07034_),
    .X(_08335_));
 sky130_fd_sc_hd__o21ai_4 _24993_ (.A1(_08332_),
    .A2(_08334_),
    .B1(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__xnor2_4 _24994_ (.A(_08331_),
    .B(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__buf_6 _24995_ (.A(_14353_),
    .X(_08338_));
 sky130_fd_sc_hd__o21a_2 _24996_ (.A1(_08338_),
    .A2(_08201_),
    .B1(_08204_),
    .X(_08339_));
 sky130_fd_sc_hd__a22o_1 _24997_ (.A1(_05955_),
    .A2(_06287_),
    .B1(_08199_),
    .B2(_07648_),
    .X(_08340_));
 sky130_fd_sc_hd__nand3_4 _24998_ (.A(_14037_),
    .B(_14042_),
    .C(_06154_),
    .Y(_08341_));
 sky130_fd_sc_hd__clkbuf_4 _24999_ (.A(_06583_),
    .X(_08342_));
 sky130_fd_sc_hd__or2b_1 _25000_ (.A(_08341_),
    .B_N(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__o2bb2ai_1 _25001_ (.A1_N(_08340_),
    .A2_N(_08343_),
    .B1(_14048_),
    .B2(_14340_),
    .Y(_08344_));
 sky130_fd_sc_hd__o2111ai_4 _25002_ (.A1(_14346_),
    .A2(_08341_),
    .B1(_05441_),
    .C1(_06577_),
    .D1(_08340_),
    .Y(_08345_));
 sky130_fd_sc_hd__nand2_4 _25003_ (.A(_08344_),
    .B(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__xnor2_4 _25004_ (.A(_08339_),
    .B(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__xnor2_4 _25005_ (.A(_08337_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__nor2_1 _25006_ (.A(_08212_),
    .B(_08218_),
    .Y(_08349_));
 sky130_fd_sc_hd__o21bai_4 _25007_ (.A1(_08211_),
    .A2(_08219_),
    .B1_N(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__o21a_4 _25008_ (.A1(_14374_),
    .A2(_08214_),
    .B1(_08217_),
    .X(_08351_));
 sky130_fd_sc_hd__a2bb2oi_4 _25009_ (.A1_N(_07668_),
    .A2_N(_08263_),
    .B1(_08262_),
    .B2(_08265_),
    .Y(_08352_));
 sky130_fd_sc_hd__and2_2 _25010_ (.A(_06355_),
    .B(_07650_),
    .X(_08353_));
 sky130_fd_sc_hd__buf_4 _25011_ (.A(_06485_),
    .X(_08354_));
 sky130_fd_sc_hd__buf_4 _25012_ (.A(_06070_),
    .X(_08355_));
 sky130_fd_sc_hd__nand3_4 _25013_ (.A(_08354_),
    .B(_08355_),
    .C(_05699_),
    .Y(_08356_));
 sky130_fd_sc_hd__buf_4 _25014_ (.A(_14026_),
    .X(_08357_));
 sky130_fd_sc_hd__a22o_2 _25015_ (.A1(_06349_),
    .A2(_05768_),
    .B1(_08357_),
    .B2(_06018_),
    .X(_08358_));
 sky130_fd_sc_hd__o21ai_4 _25016_ (.A1(_14366_),
    .A2(_08356_),
    .B1(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__xor2_4 _25017_ (.A(_08353_),
    .B(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__xnor2_4 _25018_ (.A(_08352_),
    .B(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__xor2_4 _25019_ (.A(_08351_),
    .B(_08361_),
    .X(_08362_));
 sky130_fd_sc_hd__xnor2_2 _25020_ (.A(_08350_),
    .B(_08362_),
    .Y(_08363_));
 sky130_fd_sc_hd__xor2_4 _25021_ (.A(_08348_),
    .B(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__nor2_4 _25022_ (.A(_08329_),
    .B(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__nand2_1 _25023_ (.A(_08364_),
    .B(_08329_),
    .Y(_08366_));
 sky130_fd_sc_hd__nor3b_4 _25024_ (.A(_08327_),
    .B(_08365_),
    .C_N(_08366_),
    .Y(_08367_));
 sky130_vsdinv _25025_ (.A(_08365_),
    .Y(_08368_));
 sky130_vsdinv _25026_ (.A(_08327_),
    .Y(_08369_));
 sky130_fd_sc_hd__a21oi_1 _25027_ (.A1(_08368_),
    .A2(_08366_),
    .B1(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__nor2_2 _25028_ (.A(_08367_),
    .B(_08370_),
    .Y(_08371_));
 sky130_vsdinv _25029_ (.A(_08371_),
    .Y(_08372_));
 sky130_fd_sc_hd__and2_2 _25030_ (.A(_07358_),
    .B(_05033_),
    .X(_08373_));
 sky130_fd_sc_hd__buf_4 _25031_ (.A(\pcpi_mul.rs2[29] ),
    .X(_08374_));
 sky130_fd_sc_hd__buf_4 _25032_ (.A(_13976_),
    .X(_08375_));
 sky130_fd_sc_hd__nand3_4 _25033_ (.A(_08374_),
    .B(_08375_),
    .C(_04974_),
    .Y(_08376_));
 sky130_fd_sc_hd__a22o_1 _25034_ (.A1(_07961_),
    .A2(_04898_),
    .B1(_13977_),
    .B2(_04957_),
    .X(_08377_));
 sky130_fd_sc_hd__o21ai_2 _25035_ (.A1(_14434_),
    .A2(_08376_),
    .B1(_08377_),
    .Y(_08378_));
 sky130_fd_sc_hd__xnor2_2 _25036_ (.A(_08373_),
    .B(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand3b_4 _25037_ (.A_N(_08246_),
    .B(_07945_),
    .C(_04908_),
    .Y(_08380_));
 sky130_fd_sc_hd__and2_1 _25038_ (.A(\pcpi_mul.rs2[30] ),
    .B(_04968_),
    .X(_08381_));
 sky130_fd_sc_hd__nand2_4 _25039_ (.A(\pcpi_mul.rs2[31] ),
    .B(_14447_),
    .Y(_08382_));
 sky130_fd_sc_hd__clkbuf_2 _25040_ (.A(\pcpi_mul.rs2[32] ),
    .X(_08383_));
 sky130_fd_sc_hd__nand2_2 _25041_ (.A(_14451_),
    .B(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__xor2_4 _25042_ (.A(_08382_),
    .B(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__xnor2_2 _25043_ (.A(_08381_),
    .B(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__xnor2_1 _25044_ (.A(_08380_),
    .B(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__xor2_1 _25045_ (.A(_08379_),
    .B(_08387_),
    .X(_08388_));
 sky130_fd_sc_hd__or2_1 _25046_ (.A(_08248_),
    .B(_08253_),
    .X(_08389_));
 sky130_fd_sc_hd__nand2_1 _25047_ (.A(_08388_),
    .B(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__or2b_2 _25048_ (.A(_08387_),
    .B_N(_08379_),
    .X(_08391_));
 sky130_fd_sc_hd__or2b_1 _25049_ (.A(_08379_),
    .B_N(_08387_),
    .X(_08392_));
 sky130_fd_sc_hd__nand3b_1 _25050_ (.A_N(_08389_),
    .B(_08391_),
    .C(_08392_),
    .Y(_08393_));
 sky130_fd_sc_hd__nand2_1 _25051_ (.A(_08390_),
    .B(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__o21a_1 _25052_ (.A1(_14423_),
    .A2(_08237_),
    .B1(_08240_),
    .X(_08395_));
 sky130_fd_sc_hd__buf_6 _25053_ (.A(_13971_),
    .X(_08396_));
 sky130_fd_sc_hd__buf_6 _25054_ (.A(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__nand3b_1 _25055_ (.A_N(_08250_),
    .B(_08397_),
    .C(_04891_),
    .Y(_08398_));
 sky130_fd_sc_hd__o31a_2 _25056_ (.A1(_13982_),
    .A2(_14434_),
    .A3(_08252_),
    .B1(_08398_),
    .X(_08399_));
 sky130_fd_sc_hd__buf_6 _25057_ (.A(_06887_),
    .X(_08400_));
 sky130_fd_sc_hd__nand2_2 _25058_ (.A(_08400_),
    .B(_05229_),
    .Y(_08401_));
 sky130_fd_sc_hd__buf_2 _25059_ (.A(_13984_),
    .X(_08402_));
 sky130_fd_sc_hd__or4_4 _25060_ (.A(_08402_),
    .B(_13989_),
    .C(_14416_),
    .D(_14421_),
    .X(_08403_));
 sky130_fd_sc_hd__clkbuf_4 _25061_ (.A(_07264_),
    .X(_08404_));
 sky130_fd_sc_hd__clkbuf_4 _25062_ (.A(_07265_),
    .X(_08405_));
 sky130_fd_sc_hd__a22o_1 _25063_ (.A1(_08404_),
    .A2(_05041_),
    .B1(_08405_),
    .B2(_05101_),
    .X(_08406_));
 sky130_fd_sc_hd__nand2_2 _25064_ (.A(_08403_),
    .B(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__xnor2_2 _25065_ (.A(_08401_),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__xnor2_2 _25066_ (.A(_08399_),
    .B(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__xor2_2 _25067_ (.A(_08395_),
    .B(_08409_),
    .X(_08410_));
 sky130_fd_sc_hd__xnor2_1 _25068_ (.A(_08394_),
    .B(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__or2b_1 _25069_ (.A(_08243_),
    .B_N(_08255_),
    .X(_08412_));
 sky130_fd_sc_hd__o21ai_1 _25070_ (.A1(_08245_),
    .A2(_08254_),
    .B1(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__and2_1 _25071_ (.A(_08411_),
    .B(_08413_),
    .X(_08414_));
 sky130_vsdinv _25072_ (.A(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__or2_4 _25073_ (.A(_08413_),
    .B(_08411_),
    .X(_08416_));
 sky130_fd_sc_hd__nor2_1 _25074_ (.A(_08268_),
    .B(_08275_),
    .Y(_08417_));
 sky130_fd_sc_hd__o21bai_4 _25075_ (.A1(_08267_),
    .A2(_08276_),
    .B1_N(_08417_),
    .Y(_08418_));
 sky130_fd_sc_hd__a21o_1 _25076_ (.A1(_07957_),
    .A2(_07959_),
    .B1(_08242_),
    .X(_08419_));
 sky130_fd_sc_hd__o21ai_4 _25077_ (.A1(_08235_),
    .A2(_08241_),
    .B1(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__and2_2 _25078_ (.A(_06346_),
    .B(_05611_),
    .X(_08421_));
 sky130_fd_sc_hd__buf_6 _25079_ (.A(_06895_),
    .X(_08422_));
 sky130_fd_sc_hd__buf_6 _25080_ (.A(_14015_),
    .X(_08423_));
 sky130_fd_sc_hd__nand3_4 _25081_ (.A(_08422_),
    .B(_08423_),
    .C(_05597_),
    .Y(_08424_));
 sky130_fd_sc_hd__buf_6 _25082_ (.A(_06322_),
    .X(_08425_));
 sky130_fd_sc_hd__buf_4 _25083_ (.A(_06185_),
    .X(_08426_));
 sky130_fd_sc_hd__a22o_2 _25084_ (.A1(_08425_),
    .A2(_05505_),
    .B1(_08426_),
    .B2(_06161_),
    .X(_08427_));
 sky130_fd_sc_hd__o21ai_4 _25085_ (.A1(_14385_),
    .A2(_08424_),
    .B1(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__xor2_4 _25086_ (.A(_08421_),
    .B(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__o21a_2 _25087_ (.A1(_14406_),
    .A2(_08271_),
    .B1(_08274_),
    .X(_08430_));
 sky130_fd_sc_hd__buf_4 _25088_ (.A(_06744_),
    .X(_08431_));
 sky130_fd_sc_hd__buf_6 _25089_ (.A(_06646_),
    .X(_08432_));
 sky130_fd_sc_hd__a22o_1 _25090_ (.A1(_08431_),
    .A2(_05237_),
    .B1(_08432_),
    .B2(_05614_),
    .X(_08433_));
 sky130_fd_sc_hd__nand3_4 _25091_ (.A(_07246_),
    .B(_06647_),
    .C(_05516_),
    .Y(_08434_));
 sky130_fd_sc_hd__or2b_1 _25092_ (.A(_08434_),
    .B_N(_05311_),
    .X(_08435_));
 sky130_fd_sc_hd__o2bb2ai_1 _25093_ (.A1_N(_08433_),
    .A2_N(_08435_),
    .B1(_07123_),
    .B2(_14395_),
    .Y(_08436_));
 sky130_fd_sc_hd__o2111ai_4 _25094_ (.A1(_05874_),
    .A2(_08434_),
    .B1(_06471_),
    .C1(_05414_),
    .D1(_08433_),
    .Y(_08437_));
 sky130_fd_sc_hd__nand2_4 _25095_ (.A(_08436_),
    .B(_08437_),
    .Y(_08438_));
 sky130_fd_sc_hd__xnor2_4 _25096_ (.A(_08430_),
    .B(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__xor2_4 _25097_ (.A(_08429_),
    .B(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__xnor2_4 _25098_ (.A(_08420_),
    .B(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__xnor2_4 _25099_ (.A(_08418_),
    .B(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__a21o_1 _25100_ (.A1(_08415_),
    .A2(_08416_),
    .B1(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__nand3b_4 _25101_ (.A_N(_08414_),
    .B(_08442_),
    .C(_08416_),
    .Y(_08444_));
 sky130_fd_sc_hd__a21boi_1 _25102_ (.A1(_08257_),
    .A2(_08281_),
    .B1_N(_08258_),
    .Y(_08445_));
 sky130_vsdinv _25103_ (.A(_08445_),
    .Y(_08446_));
 sky130_fd_sc_hd__a21oi_4 _25104_ (.A1(_08443_),
    .A2(_08444_),
    .B1(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__nand3_1 _25105_ (.A(_08443_),
    .B(_08444_),
    .C(_08446_),
    .Y(_08448_));
 sky130_vsdinv _25106_ (.A(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__nor3_4 _25107_ (.A(_08372_),
    .B(_08447_),
    .C(_08449_),
    .Y(_08450_));
 sky130_vsdinv _25108_ (.A(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__o21bai_4 _25109_ (.A1(_08447_),
    .A2(_08449_),
    .B1_N(_08371_),
    .Y(_08452_));
 sky130_fd_sc_hd__o21a_1 _25110_ (.A1(_08231_),
    .A2(_08286_),
    .B1(_08284_),
    .X(_08453_));
 sky130_vsdinv _25111_ (.A(_08453_),
    .Y(_08454_));
 sky130_fd_sc_hd__a21oi_4 _25112_ (.A1(_08451_),
    .A2(_08452_),
    .B1(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__nand3_4 _25113_ (.A(_08454_),
    .B(_08451_),
    .C(_08452_),
    .Y(_08456_));
 sky130_vsdinv _25114_ (.A(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__a21boi_4 _25115_ (.A1(_08180_),
    .A2(_08154_),
    .B1_N(_08155_),
    .Y(_08458_));
 sky130_fd_sc_hd__nor2_1 _25116_ (.A(_08141_),
    .B(_08146_),
    .Y(_08459_));
 sky130_fd_sc_hd__o21ba_1 _25117_ (.A1(_08140_),
    .A2(_08147_),
    .B1_N(_08459_),
    .X(_08460_));
 sky130_vsdinv _25118_ (.A(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__or2b_1 _25119_ (.A(_08206_),
    .B_N(_08197_),
    .X(_08462_));
 sky130_fd_sc_hd__o21ai_4 _25120_ (.A1(_08205_),
    .A2(_08198_),
    .B1(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__buf_8 _25121_ (.A(_14315_),
    .X(_08464_));
 sky130_fd_sc_hd__a2bb2oi_4 _25122_ (.A1_N(_08464_),
    .A2_N(_08143_),
    .B1(_08142_),
    .B2(_08144_),
    .Y(_08465_));
 sky130_fd_sc_hd__a2bb2oi_4 _25123_ (.A1_N(_07214_),
    .A2_N(_08194_),
    .B1(_08193_),
    .B2(_08195_),
    .Y(_08466_));
 sky130_fd_sc_hd__and2_2 _25124_ (.A(_04997_),
    .B(_07216_),
    .X(_08467_));
 sky130_fd_sc_hd__nand3_4 _25125_ (.A(_05126_),
    .B(_05064_),
    .C(_07038_),
    .Y(_08468_));
 sky130_fd_sc_hd__a22o_2 _25126_ (.A1(_05131_),
    .A2(_06956_),
    .B1(_05064_),
    .B2(_07786_),
    .X(_08469_));
 sky130_fd_sc_hd__o21ai_4 _25127_ (.A1(_14308_),
    .A2(_08468_),
    .B1(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__xor2_4 _25128_ (.A(_08467_),
    .B(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__xnor2_4 _25129_ (.A(_08466_),
    .B(_08471_),
    .Y(_08472_));
 sky130_fd_sc_hd__xor2_4 _25130_ (.A(_08465_),
    .B(_08472_),
    .X(_08473_));
 sky130_fd_sc_hd__xnor2_4 _25131_ (.A(_08463_),
    .B(_08473_),
    .Y(_08474_));
 sky130_fd_sc_hd__xor2_4 _25132_ (.A(_08461_),
    .B(_08474_),
    .X(_08475_));
 sky130_fd_sc_hd__a21oi_2 _25133_ (.A1(_08139_),
    .A2(_08148_),
    .B1(_08150_),
    .Y(_08476_));
 sky130_fd_sc_hd__nand2_2 _25134_ (.A(_08475_),
    .B(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__nor2_2 _25135_ (.A(_08476_),
    .B(_08475_),
    .Y(_08478_));
 sky130_vsdinv _25136_ (.A(_08478_),
    .Y(_08479_));
 sky130_fd_sc_hd__buf_2 _25137_ (.A(_08165_),
    .X(_08480_));
 sky130_fd_sc_hd__buf_2 _25138_ (.A(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__buf_4 _25139_ (.A(_08481_),
    .X(_08482_));
 sky130_fd_sc_hd__nor3_4 _25140_ (.A(_14088_),
    .B(_14294_),
    .C(_08167_),
    .Y(_08483_));
 sky130_fd_sc_hd__a41oi_4 _25141_ (.A1(_05299_),
    .A2(_04880_),
    .A3(_08482_),
    .A4(_08158_),
    .B1(_08483_),
    .Y(_08484_));
 sky130_fd_sc_hd__nor2_1 _25142_ (.A(_08169_),
    .B(_08176_),
    .Y(_08485_));
 sky130_fd_sc_hd__o21bai_4 _25143_ (.A1(_08168_),
    .A2(_08177_),
    .B1_N(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__buf_2 _25144_ (.A(\pcpi_mul.rs1[29] ),
    .X(_08487_));
 sky130_fd_sc_hd__clkbuf_4 _25145_ (.A(_08487_),
    .X(_08488_));
 sky130_fd_sc_hd__buf_2 _25146_ (.A(_08488_),
    .X(_08489_));
 sky130_fd_sc_hd__and2_2 _25147_ (.A(_14084_),
    .B(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__nand2_2 _25148_ (.A(_04885_),
    .B(_08480_),
    .Y(_08491_));
 sky130_fd_sc_hd__buf_2 _25149_ (.A(_08171_),
    .X(_08492_));
 sky130_fd_sc_hd__nand2_2 _25150_ (.A(_04877_),
    .B(_08492_),
    .Y(_08493_));
 sky130_fd_sc_hd__xnor2_4 _25151_ (.A(_08491_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__xor2_4 _25152_ (.A(_08490_),
    .B(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__o21a_2 _25153_ (.A1(_08172_),
    .A2(_08175_),
    .B1(_08173_),
    .X(_08496_));
 sky130_fd_sc_hd__and2_1 _25154_ (.A(_12777_),
    .B(_05045_),
    .X(_08497_));
 sky130_fd_sc_hd__buf_6 _25155_ (.A(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__or4_4 _25156_ (.A(_14074_),
    .B(_14077_),
    .C(_14290_),
    .D(_14296_),
    .X(_08499_));
 sky130_fd_sc_hd__a22o_2 _25157_ (.A1(_05117_),
    .A2(_07485_),
    .B1(_05515_),
    .B2(_07585_),
    .X(_08500_));
 sky130_fd_sc_hd__nand2_2 _25158_ (.A(_08499_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__xor2_4 _25159_ (.A(_08498_),
    .B(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__xnor2_4 _25160_ (.A(_08496_),
    .B(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__xor2_4 _25161_ (.A(_08495_),
    .B(_08503_),
    .X(_08504_));
 sky130_fd_sc_hd__xnor2_4 _25162_ (.A(_08486_),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__xor2_4 _25163_ (.A(_08484_),
    .B(_08505_),
    .X(_08506_));
 sky130_fd_sc_hd__a21oi_4 _25164_ (.A1(_08477_),
    .A2(_08479_),
    .B1(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__and3_2 _25165_ (.A(_08506_),
    .B(_08479_),
    .C(_08477_),
    .X(_08508_));
 sky130_fd_sc_hd__and2_1 _25166_ (.A(_08230_),
    .B(_08226_),
    .X(_08509_));
 sky130_fd_sc_hd__o21a_2 _25167_ (.A1(_08507_),
    .A2(_08508_),
    .B1(_08509_),
    .X(_08510_));
 sky130_fd_sc_hd__a211oi_4 _25168_ (.A1(_08226_),
    .A2(_08230_),
    .B1(_08507_),
    .C1(_08508_),
    .Y(_08511_));
 sky130_fd_sc_hd__nor3_4 _25169_ (.A(_08458_),
    .B(_08510_),
    .C(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__o21a_1 _25170_ (.A1(_08510_),
    .A2(_08511_),
    .B1(_08458_),
    .X(_08513_));
 sky130_fd_sc_hd__nor2_4 _25171_ (.A(_08512_),
    .B(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__o21bai_4 _25172_ (.A1(_08455_),
    .A2(_08457_),
    .B1_N(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__nand3b_4 _25173_ (.A_N(_08455_),
    .B(_08514_),
    .C(_08456_),
    .Y(_08516_));
 sky130_fd_sc_hd__nand2_1 _25174_ (.A(_08515_),
    .B(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__a21boi_2 _25175_ (.A1(_08192_),
    .A2(_08292_),
    .B1_N(_08291_),
    .Y(_08518_));
 sky130_fd_sc_hd__nand2_2 _25176_ (.A(_08517_),
    .B(_08518_),
    .Y(_08519_));
 sky130_vsdinv _25177_ (.A(_08518_),
    .Y(_08520_));
 sky130_fd_sc_hd__nand3_4 _25178_ (.A(_08520_),
    .B(_08515_),
    .C(_08516_),
    .Y(_08521_));
 sky130_fd_sc_hd__nand2_1 _25179_ (.A(_08178_),
    .B(_08162_),
    .Y(_08522_));
 sky130_fd_sc_hd__o21a_4 _25180_ (.A1(_08160_),
    .A2(_08179_),
    .B1(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__a21o_2 _25181_ (.A1(_08190_),
    .A2(_08186_),
    .B1(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__nand3_4 _25182_ (.A(_08190_),
    .B(_08186_),
    .C(_08523_),
    .Y(_08525_));
 sky130_fd_sc_hd__buf_6 _25183_ (.A(_12805_),
    .X(_08526_));
 sky130_fd_sc_hd__buf_2 _25184_ (.A(_08526_),
    .X(_08527_));
 sky130_fd_sc_hd__clkbuf_4 _25185_ (.A(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__clkbuf_4 _25186_ (.A(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__a21oi_2 _25187_ (.A1(_08524_),
    .A2(_08525_),
    .B1(net420),
    .Y(_08530_));
 sky130_fd_sc_hd__nand3_4 _25188_ (.A(_08524_),
    .B(net420),
    .C(_08525_),
    .Y(_08531_));
 sky130_fd_sc_hd__and2b_1 _25189_ (.A_N(_08530_),
    .B(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__a21oi_1 _25190_ (.A1(_08519_),
    .A2(_08521_),
    .B1(_08532_),
    .Y(_08533_));
 sky130_fd_sc_hd__nand3_4 _25191_ (.A(_08519_),
    .B(_08532_),
    .C(_08521_),
    .Y(_08534_));
 sky130_vsdinv _25192_ (.A(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__a21o_1 _25193_ (.A1(_08304_),
    .A2(_08302_),
    .B1(_08298_),
    .X(_08536_));
 sky130_fd_sc_hd__o21bai_2 _25194_ (.A1(_08533_),
    .A2(_08535_),
    .B1_N(_08536_),
    .Y(_08537_));
 sky130_vsdinv _25195_ (.A(_08531_),
    .Y(_08538_));
 sky130_fd_sc_hd__o2bb2ai_2 _25196_ (.A1_N(_08521_),
    .A2_N(_08519_),
    .B1(_08538_),
    .B2(_08530_),
    .Y(_08539_));
 sky130_fd_sc_hd__nand3_4 _25197_ (.A(_08539_),
    .B(_08534_),
    .C(_08536_),
    .Y(_08540_));
 sky130_fd_sc_hd__and2_1 _25198_ (.A(_08301_),
    .B(_08300_),
    .X(_08541_));
 sky130_fd_sc_hd__a21o_1 _25199_ (.A1(_08537_),
    .A2(_08540_),
    .B1(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__nand3_4 _25200_ (.A(_08537_),
    .B(_08540_),
    .C(_08541_),
    .Y(_08543_));
 sky130_fd_sc_hd__nand2_2 _25201_ (.A(_08313_),
    .B(_08310_),
    .Y(_08544_));
 sky130_fd_sc_hd__a21o_1 _25202_ (.A1(_08542_),
    .A2(_08543_),
    .B1(_08544_),
    .X(_08545_));
 sky130_fd_sc_hd__nand3_4 _25203_ (.A(_08542_),
    .B(_08543_),
    .C(_08544_),
    .Y(_08546_));
 sky130_fd_sc_hd__nand2_4 _25204_ (.A(_08545_),
    .B(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__o21bai_1 _25205_ (.A1(_08319_),
    .A2(_08320_),
    .B1_N(_08316_),
    .Y(_08548_));
 sky130_fd_sc_hd__nand3_2 _25206_ (.A(_08312_),
    .B(_08313_),
    .C(_08316_),
    .Y(_08549_));
 sky130_fd_sc_hd__nand2_1 _25207_ (.A(_08548_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__nor2_1 _25208_ (.A(_08130_),
    .B(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__nand2_2 _25209_ (.A(_08551_),
    .B(_08132_),
    .Y(_08552_));
 sky130_fd_sc_hd__nor2_4 _25210_ (.A(_07738_),
    .B(_08552_),
    .Y(_08553_));
 sky130_fd_sc_hd__nand3_4 _25211_ (.A(_05867_),
    .B(_08553_),
    .C(_07000_),
    .Y(_08554_));
 sky130_fd_sc_hd__nand2_4 _25212_ (.A(_07005_),
    .B(_08553_),
    .Y(_08555_));
 sky130_fd_sc_hd__a21oi_1 _25213_ (.A1(_07720_),
    .A2(_07723_),
    .B1(_07727_),
    .Y(_08556_));
 sky130_fd_sc_hd__nor3_2 _25214_ (.A(_08556_),
    .B(_07931_),
    .C(_07933_),
    .Y(_08557_));
 sky130_fd_sc_hd__nor2_1 _25215_ (.A(_08133_),
    .B(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__nand2_1 _25216_ (.A(_07734_),
    .B(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__nor2_1 _25217_ (.A(_08323_),
    .B(_08324_),
    .Y(_08560_));
 sky130_fd_sc_hd__nand2_1 _25218_ (.A(_08322_),
    .B(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__nor2_2 _25219_ (.A(_08559_),
    .B(_08561_),
    .Y(_08562_));
 sky130_fd_sc_hd__nand3_1 _25220_ (.A(_08322_),
    .B(_08560_),
    .C(_08134_),
    .Y(_08563_));
 sky130_fd_sc_hd__nand2_1 _25221_ (.A(_08324_),
    .B(_08548_),
    .Y(_08564_));
 sky130_fd_sc_hd__nand3_2 _25222_ (.A(_08563_),
    .B(_08549_),
    .C(_08564_),
    .Y(_08565_));
 sky130_fd_sc_hd__a21oi_4 _25223_ (.A1(_08562_),
    .A2(_07744_),
    .B1(_08565_),
    .Y(_08566_));
 sky130_fd_sc_hd__nand3_4 _25224_ (.A(_08554_),
    .B(_08555_),
    .C(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__xnor2_1 _25225_ (.A(_08547_),
    .B(_08567_),
    .Y(_02651_));
 sky130_fd_sc_hd__nand2_2 _25226_ (.A(_08473_),
    .B(_08463_),
    .Y(_08568_));
 sky130_fd_sc_hd__or2b_2 _25227_ (.A(_08474_),
    .B_N(_08461_),
    .X(_08569_));
 sky130_fd_sc_hd__nor2_1 _25228_ (.A(_08466_),
    .B(_08471_),
    .Y(_08570_));
 sky130_fd_sc_hd__o21ba_1 _25229_ (.A1(_08465_),
    .A2(_08472_),
    .B1_N(_08570_),
    .X(_08571_));
 sky130_fd_sc_hd__or2b_1 _25230_ (.A(_08347_),
    .B_N(_08337_),
    .X(_08572_));
 sky130_fd_sc_hd__o21ai_2 _25231_ (.A1(_08346_),
    .A2(_08339_),
    .B1(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__a2bb2oi_4 _25232_ (.A1_N(_14311_),
    .A2_N(_08468_),
    .B1(_08467_),
    .B2(_08469_),
    .Y(_08574_));
 sky130_fd_sc_hd__a2bb2oi_4 _25233_ (.A1_N(_08332_),
    .A2_N(_08334_),
    .B1(_08331_),
    .B2(_08335_),
    .Y(_08575_));
 sky130_fd_sc_hd__nand2_4 _25234_ (.A(_04999_),
    .B(_07769_),
    .Y(_08576_));
 sky130_fd_sc_hd__or4_4 _25235_ (.A(_14063_),
    .B(_14067_),
    .C(_14303_),
    .D(_14308_),
    .X(_08577_));
 sky130_fd_sc_hd__a22o_1 _25236_ (.A1(_05132_),
    .A2(_07044_),
    .B1(_05164_),
    .B2(_07477_),
    .X(_08578_));
 sky130_fd_sc_hd__nand2_2 _25237_ (.A(_08577_),
    .B(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__xnor2_4 _25238_ (.A(_08576_),
    .B(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__xnor2_4 _25239_ (.A(_08575_),
    .B(_08580_),
    .Y(_08581_));
 sky130_fd_sc_hd__xor2_4 _25240_ (.A(_08574_),
    .B(_08581_),
    .X(_08582_));
 sky130_fd_sc_hd__xnor2_2 _25241_ (.A(_08573_),
    .B(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__xnor2_2 _25242_ (.A(_08571_),
    .B(_08583_),
    .Y(_08584_));
 sky130_fd_sc_hd__a21o_1 _25243_ (.A1(_08568_),
    .A2(_08569_),
    .B1(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__nand3_4 _25244_ (.A(_08584_),
    .B(_08568_),
    .C(_08569_),
    .Y(_08586_));
 sky130_fd_sc_hd__nand2_1 _25245_ (.A(_08585_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__clkbuf_4 _25246_ (.A(_08492_),
    .X(_08588_));
 sky130_fd_sc_hd__buf_4 _25247_ (.A(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__nor3_4 _25248_ (.A(_14088_),
    .B(_14287_),
    .C(_08494_),
    .Y(_08590_));
 sky130_fd_sc_hd__a41oi_4 _25249_ (.A1(_05299_),
    .A2(_04880_),
    .A3(_08589_),
    .A4(_08482_),
    .B1(_08590_),
    .Y(_08591_));
 sky130_fd_sc_hd__nor2_1 _25250_ (.A(_08496_),
    .B(_08502_),
    .Y(_08592_));
 sky130_fd_sc_hd__o21bai_4 _25251_ (.A1(_08495_),
    .A2(_08503_),
    .B1_N(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__and2_2 _25252_ (.A(_14084_),
    .B(_08481_),
    .X(_08594_));
 sky130_fd_sc_hd__clkbuf_4 _25253_ (.A(_08171_),
    .X(_08595_));
 sky130_fd_sc_hd__buf_4 _25254_ (.A(_08595_),
    .X(_08596_));
 sky130_fd_sc_hd__nand2_2 _25255_ (.A(_04885_),
    .B(_08596_),
    .Y(_08597_));
 sky130_fd_sc_hd__nand2_8 _25256_ (.A(_12776_),
    .B(\pcpi_mul.rs2[1] ),
    .Y(_08598_));
 sky130_fd_sc_hd__xnor2_4 _25257_ (.A(_08597_),
    .B(_08598_),
    .Y(_08599_));
 sky130_fd_sc_hd__xor2_4 _25258_ (.A(_08594_),
    .B(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__buf_8 _25259_ (.A(_08498_),
    .X(_08601_));
 sky130_fd_sc_hd__a21boi_4 _25260_ (.A1(_08500_),
    .A2(_08601_),
    .B1_N(_08499_),
    .Y(_08602_));
 sky130_fd_sc_hd__or4_4 _25261_ (.A(_14075_),
    .B(_14077_),
    .C(_08084_),
    .D(_14291_),
    .X(_08603_));
 sky130_fd_sc_hd__clkbuf_4 _25262_ (.A(_05515_),
    .X(_08604_));
 sky130_fd_sc_hd__a22o_2 _25263_ (.A1(_06159_),
    .A2(_07778_),
    .B1(_08604_),
    .B2(_08488_),
    .X(_08605_));
 sky130_fd_sc_hd__nand2_2 _25264_ (.A(_08603_),
    .B(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__xor2_4 _25265_ (.A(_08601_),
    .B(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__xnor2_4 _25266_ (.A(_08602_),
    .B(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__xor2_4 _25267_ (.A(_08600_),
    .B(_08608_),
    .X(_08609_));
 sky130_fd_sc_hd__xnor2_4 _25268_ (.A(_08593_),
    .B(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__xor2_4 _25269_ (.A(_08591_),
    .B(_08610_),
    .X(_08611_));
 sky130_vsdinv _25270_ (.A(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__nand2_2 _25271_ (.A(_08587_),
    .B(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__nand3_4 _25272_ (.A(_08585_),
    .B(_08586_),
    .C(_08611_),
    .Y(_08614_));
 sky130_fd_sc_hd__a21o_2 _25273_ (.A1(_08366_),
    .A2(_08369_),
    .B1(_08365_),
    .X(_08615_));
 sky130_fd_sc_hd__a21o_2 _25274_ (.A1(_08613_),
    .A2(_08614_),
    .B1(_08615_),
    .X(_08616_));
 sky130_fd_sc_hd__nand3_4 _25275_ (.A(_08613_),
    .B(_08615_),
    .C(_08614_),
    .Y(_08617_));
 sky130_fd_sc_hd__a21oi_1 _25276_ (.A1(_08506_),
    .A2(_08477_),
    .B1(_08478_),
    .Y(_08618_));
 sky130_fd_sc_hd__a21boi_4 _25277_ (.A1(_08616_),
    .A2(_08617_),
    .B1_N(_08618_),
    .Y(_08619_));
 sky130_fd_sc_hd__o211a_4 _25278_ (.A1(_08478_),
    .A2(_08508_),
    .B1(_08617_),
    .C1(_08616_),
    .X(_08620_));
 sky130_fd_sc_hd__nor2_2 _25279_ (.A(_08619_),
    .B(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__a21bo_2 _25280_ (.A1(_08410_),
    .A2(_08390_),
    .B1_N(_08393_),
    .X(_08622_));
 sky130_fd_sc_hd__o21a_2 _25281_ (.A1(_08401_),
    .A2(_08407_),
    .B1(_08403_),
    .X(_08623_));
 sky130_fd_sc_hd__a2bb2oi_4 _25282_ (.A1_N(_14435_),
    .A2_N(_08376_),
    .B1(_08373_),
    .B2(_08377_),
    .Y(_08624_));
 sky130_fd_sc_hd__nand2_4 _25283_ (.A(_06888_),
    .B(_05301_),
    .Y(_08625_));
 sky130_fd_sc_hd__or4_4 _25284_ (.A(_13985_),
    .B(_13990_),
    .C(_05998_),
    .D(_14417_),
    .X(_08626_));
 sky130_fd_sc_hd__buf_4 _25285_ (.A(_07264_),
    .X(_08627_));
 sky130_fd_sc_hd__buf_4 _25286_ (.A(_07265_),
    .X(_08628_));
 sky130_fd_sc_hd__a22o_1 _25287_ (.A1(_08627_),
    .A2(_05819_),
    .B1(_08628_),
    .B2(_05228_),
    .X(_08629_));
 sky130_fd_sc_hd__nand2_2 _25288_ (.A(_08626_),
    .B(_08629_),
    .Y(_08630_));
 sky130_fd_sc_hd__xnor2_4 _25289_ (.A(_08625_),
    .B(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__xnor2_4 _25290_ (.A(_08624_),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__xor2_4 _25291_ (.A(_08623_),
    .B(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__clkbuf_2 _25292_ (.A(\pcpi_mul.rs2[27] ),
    .X(_08634_));
 sky130_fd_sc_hd__and2_2 _25293_ (.A(_08634_),
    .B(_05092_),
    .X(_08635_));
 sky130_fd_sc_hd__clkbuf_4 _25294_ (.A(_13971_),
    .X(_08636_));
 sky130_fd_sc_hd__buf_6 _25295_ (.A(_13977_),
    .X(_08637_));
 sky130_fd_sc_hd__nand3_4 _25296_ (.A(_08636_),
    .B(_08637_),
    .C(_04928_),
    .Y(_08638_));
 sky130_fd_sc_hd__a22o_2 _25297_ (.A1(_07961_),
    .A2(_04957_),
    .B1(_08375_),
    .B2(_05039_),
    .X(_08639_));
 sky130_fd_sc_hd__o21ai_4 _25298_ (.A1(_05247_),
    .A2(_08638_),
    .B1(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__xor2_4 _25299_ (.A(_08635_),
    .B(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__nor3_4 _25300_ (.A(_04717_),
    .B(_12806_),
    .C(_08382_),
    .Y(_08642_));
 sky130_fd_sc_hd__a21o_2 _25301_ (.A1(_08385_),
    .A2(_08381_),
    .B1(_08642_),
    .X(_08643_));
 sky130_fd_sc_hd__clkbuf_2 _25302_ (.A(\pcpi_mul.rs2[30] ),
    .X(_08644_));
 sky130_fd_sc_hd__and2_2 _25303_ (.A(_08644_),
    .B(_04898_),
    .X(_08645_));
 sky130_fd_sc_hd__clkbuf_4 _25304_ (.A(\pcpi_mul.rs2[31] ),
    .X(_08646_));
 sky130_fd_sc_hd__nand2_2 _25305_ (.A(_08646_),
    .B(_04889_),
    .Y(_08647_));
 sky130_fd_sc_hd__and2b_1 _25306_ (.A_N(_04906_),
    .B(_08383_),
    .X(_08648_));
 sky130_fd_sc_hd__xor2_4 _25307_ (.A(_08647_),
    .B(_08648_),
    .X(_08649_));
 sky130_fd_sc_hd__xor2_4 _25308_ (.A(_08645_),
    .B(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__xor2_4 _25309_ (.A(_08643_),
    .B(_08650_),
    .X(_08651_));
 sky130_fd_sc_hd__xor2_4 _25310_ (.A(_08641_),
    .B(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__o21ai_4 _25311_ (.A1(_08380_),
    .A2(_08386_),
    .B1(_08391_),
    .Y(_08653_));
 sky130_fd_sc_hd__xnor2_2 _25312_ (.A(_08652_),
    .B(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__xnor2_2 _25313_ (.A(_08633_),
    .B(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__nor2_4 _25314_ (.A(_08622_),
    .B(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__nor2_1 _25315_ (.A(_08430_),
    .B(_08438_),
    .Y(_08657_));
 sky130_fd_sc_hd__o21ba_1 _25316_ (.A1(_08429_),
    .A2(_08439_),
    .B1_N(_08657_),
    .X(_08658_));
 sky130_fd_sc_hd__and2_2 _25317_ (.A(_08261_),
    .B(_05905_),
    .X(_08659_));
 sky130_fd_sc_hd__buf_6 _25318_ (.A(_14010_),
    .X(_08660_));
 sky130_fd_sc_hd__nand3_4 _25319_ (.A(_08660_),
    .B(_08426_),
    .C(_06161_),
    .Y(_08661_));
 sky130_fd_sc_hd__clkbuf_4 _25320_ (.A(_06322_),
    .X(_08662_));
 sky130_fd_sc_hd__a22o_2 _25321_ (.A1(_08662_),
    .A2(_05513_),
    .B1(_06896_),
    .B2(_05691_),
    .X(_08663_));
 sky130_fd_sc_hd__o21ai_4 _25322_ (.A1(_14379_),
    .A2(_08661_),
    .B1(_08663_),
    .Y(_08664_));
 sky130_fd_sc_hd__xor2_4 _25323_ (.A(_08659_),
    .B(_08664_),
    .X(_08665_));
 sky130_fd_sc_hd__o21a_2 _25324_ (.A1(_14401_),
    .A2(_08434_),
    .B1(_08437_),
    .X(_08666_));
 sky130_fd_sc_hd__buf_4 _25325_ (.A(_13998_),
    .X(_08667_));
 sky130_fd_sc_hd__clkbuf_4 _25326_ (.A(_07979_),
    .X(_08668_));
 sky130_fd_sc_hd__a22o_1 _25327_ (.A1(_08667_),
    .A2(_05614_),
    .B1(_08668_),
    .B2(_05497_),
    .X(_08669_));
 sky130_fd_sc_hd__nand3_4 _25328_ (.A(_08269_),
    .B(_07979_),
    .C(_05614_),
    .Y(_08670_));
 sky130_fd_sc_hd__or2b_1 _25329_ (.A(_08670_),
    .B_N(_05322_),
    .X(_08671_));
 sky130_fd_sc_hd__o2bb2ai_1 _25330_ (.A1_N(_08669_),
    .A2_N(_08671_),
    .B1(_07123_),
    .B2(_07668_),
    .Y(_08672_));
 sky130_fd_sc_hd__buf_6 _25331_ (.A(_06649_),
    .X(_08673_));
 sky130_fd_sc_hd__o2111ai_4 _25332_ (.A1(_05418_),
    .A2(_08670_),
    .B1(_08673_),
    .C1(_05505_),
    .D1(_08669_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand2_2 _25333_ (.A(_08672_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__xnor2_2 _25334_ (.A(_08666_),
    .B(_08675_),
    .Y(_08676_));
 sky130_fd_sc_hd__xor2_2 _25335_ (.A(_08665_),
    .B(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__nor2_1 _25336_ (.A(_08399_),
    .B(_08408_),
    .Y(_08678_));
 sky130_fd_sc_hd__o21bai_2 _25337_ (.A1(_08395_),
    .A2(_08409_),
    .B1_N(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__xnor2_1 _25338_ (.A(_08677_),
    .B(_08679_),
    .Y(_08680_));
 sky130_fd_sc_hd__xor2_1 _25339_ (.A(_08658_),
    .B(_08680_),
    .X(_08681_));
 sky130_vsdinv _25340_ (.A(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__nand2_2 _25341_ (.A(_08655_),
    .B(_08622_),
    .Y(_08683_));
 sky130_fd_sc_hd__nor3b_4 _25342_ (.A(_08656_),
    .B(_08682_),
    .C_N(_08683_),
    .Y(_08684_));
 sky130_fd_sc_hd__and2_1 _25343_ (.A(_08655_),
    .B(_08622_),
    .X(_08685_));
 sky130_fd_sc_hd__o21a_1 _25344_ (.A1(_08656_),
    .A2(_08685_),
    .B1(_08682_),
    .X(_08686_));
 sky130_fd_sc_hd__a21oi_4 _25345_ (.A1(_08416_),
    .A2(_08442_),
    .B1(_08414_),
    .Y(_08687_));
 sky130_fd_sc_hd__o21a_2 _25346_ (.A1(_08684_),
    .A2(_08686_),
    .B1(_08687_),
    .X(_08688_));
 sky130_vsdinv _25347_ (.A(_08688_),
    .Y(_08689_));
 sky130_fd_sc_hd__nor3_4 _25348_ (.A(_08687_),
    .B(_08684_),
    .C(_08686_),
    .Y(_08690_));
 sky130_vsdinv _25349_ (.A(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__xor2_2 _25350_ (.A(_08350_),
    .B(_08362_),
    .X(_08692_));
 sky130_fd_sc_hd__and2_1 _25351_ (.A(_08362_),
    .B(_08350_),
    .X(_08693_));
 sky130_fd_sc_hd__a21oi_4 _25352_ (.A1(_08692_),
    .A2(_08348_),
    .B1(_08693_),
    .Y(_08694_));
 sky130_fd_sc_hd__o21ba_1 _25353_ (.A1(_08267_),
    .A2(_08276_),
    .B1_N(_08417_),
    .X(_08695_));
 sky130_fd_sc_hd__nand2_1 _25354_ (.A(_08440_),
    .B(_08420_),
    .Y(_08696_));
 sky130_fd_sc_hd__o21a_2 _25355_ (.A1(_08695_),
    .A2(_08441_),
    .B1(_08696_),
    .X(_08697_));
 sky130_fd_sc_hd__and2_2 _25356_ (.A(_05355_),
    .B(_07198_),
    .X(_08698_));
 sky130_fd_sc_hd__buf_6 _25357_ (.A(_14320_),
    .X(_08699_));
 sky130_fd_sc_hd__nand3_4 _25358_ (.A(_05362_),
    .B(_05364_),
    .C(_07034_),
    .Y(_08700_));
 sky130_fd_sc_hd__buf_4 _25359_ (.A(_06939_),
    .X(_08701_));
 sky130_fd_sc_hd__a22o_2 _25360_ (.A1(_05362_),
    .A2(_08701_),
    .B1(_05273_),
    .B2(_07027_),
    .X(_08702_));
 sky130_fd_sc_hd__o21ai_4 _25361_ (.A1(_08699_),
    .A2(_08700_),
    .B1(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__xnor2_4 _25362_ (.A(_08698_),
    .B(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__o21a_2 _25363_ (.A1(_06293_),
    .A2(_08341_),
    .B1(_08345_),
    .X(_08705_));
 sky130_fd_sc_hd__a22o_1 _25364_ (.A1(_14037_),
    .A2(_07648_),
    .B1(_14042_),
    .B2(_06296_),
    .X(_08706_));
 sky130_fd_sc_hd__nand3_4 _25365_ (.A(_05955_),
    .B(_08199_),
    .C(_06164_),
    .Y(_08707_));
 sky130_fd_sc_hd__or2b_1 _25366_ (.A(_08707_),
    .B_N(_07746_),
    .X(_08708_));
 sky130_fd_sc_hd__o2bb2ai_1 _25367_ (.A1_N(_08706_),
    .A2_N(_08708_),
    .B1(_14047_),
    .B2(_14333_),
    .Y(_08709_));
 sky130_fd_sc_hd__buf_6 _25368_ (.A(_05532_),
    .X(_08710_));
 sky130_fd_sc_hd__o2111ai_4 _25369_ (.A1(_14339_),
    .A2(_08707_),
    .B1(_08710_),
    .C1(_06450_),
    .D1(_08706_),
    .Y(_08711_));
 sky130_fd_sc_hd__nand2_2 _25370_ (.A(_08709_),
    .B(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__xnor2_2 _25371_ (.A(_08705_),
    .B(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__xnor2_2 _25372_ (.A(_08704_),
    .B(_08713_),
    .Y(_08714_));
 sky130_vsdinv _25373_ (.A(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__nor2_1 _25374_ (.A(_08352_),
    .B(_08360_),
    .Y(_08716_));
 sky130_fd_sc_hd__o21bai_4 _25375_ (.A1(_08351_),
    .A2(_08361_),
    .B1_N(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__a2bb2oi_4 _25376_ (.A1_N(_14368_),
    .A2_N(_08356_),
    .B1(_08353_),
    .B2(_08358_),
    .Y(_08718_));
 sky130_fd_sc_hd__a2bb2oi_4 _25377_ (.A1_N(_14385_),
    .A2_N(_08424_),
    .B1(_08421_),
    .B2(_08427_),
    .Y(_08719_));
 sky130_fd_sc_hd__clkbuf_4 _25378_ (.A(_06018_),
    .X(_08720_));
 sky130_fd_sc_hd__buf_4 _25379_ (.A(_08355_),
    .X(_08721_));
 sky130_fd_sc_hd__a22o_1 _25380_ (.A1(_07294_),
    .A2(_08720_),
    .B1(_08721_),
    .B2(_05913_),
    .X(_08722_));
 sky130_fd_sc_hd__nand3_4 _25381_ (.A(_08354_),
    .B(_08355_),
    .C(_06018_),
    .Y(_08723_));
 sky130_fd_sc_hd__or2b_1 _25382_ (.A(_08723_),
    .B_N(_06030_),
    .X(_08724_));
 sky130_fd_sc_hd__o2bb2ai_1 _25383_ (.A1_N(_08722_),
    .A2_N(_08724_),
    .B1(_14032_),
    .B2(_08338_),
    .Y(_08725_));
 sky130_fd_sc_hd__o2111ai_4 _25384_ (.A1(_06034_),
    .A2(_08723_),
    .B1(net438),
    .C1(_06438_),
    .D1(_08722_),
    .Y(_08726_));
 sky130_fd_sc_hd__nand2_4 _25385_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__xnor2_4 _25386_ (.A(_08719_),
    .B(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__xor2_4 _25387_ (.A(_08718_),
    .B(_08728_),
    .X(_08729_));
 sky130_fd_sc_hd__xnor2_4 _25388_ (.A(_08717_),
    .B(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__xor2_4 _25389_ (.A(_08715_),
    .B(_08730_),
    .X(_08731_));
 sky130_fd_sc_hd__xor2_4 _25390_ (.A(_08697_),
    .B(_08731_),
    .X(_08732_));
 sky130_fd_sc_hd__xor2_4 _25391_ (.A(_08694_),
    .B(_08732_),
    .X(_08733_));
 sky130_fd_sc_hd__nand3_4 _25392_ (.A(_08689_),
    .B(_08691_),
    .C(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__o21bai_4 _25393_ (.A1(_08690_),
    .A2(_08688_),
    .B1_N(_08733_),
    .Y(_08735_));
 sky130_fd_sc_hd__o21a_1 _25394_ (.A1(_08372_),
    .A2(_08447_),
    .B1(_08448_),
    .X(_08736_));
 sky130_fd_sc_hd__a21boi_4 _25395_ (.A1(_08734_),
    .A2(_08735_),
    .B1_N(_08736_),
    .Y(_08737_));
 sky130_vsdinv _25396_ (.A(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__nand3b_4 _25397_ (.A_N(_08736_),
    .B(_08734_),
    .C(_08735_),
    .Y(_08739_));
 sky130_fd_sc_hd__nand3_4 _25398_ (.A(_08621_),
    .B(_08738_),
    .C(_08739_),
    .Y(_08740_));
 sky130_vsdinv _25399_ (.A(_08739_),
    .Y(_08741_));
 sky130_fd_sc_hd__o22ai_4 _25400_ (.A1(_08620_),
    .A2(_08619_),
    .B1(_08737_),
    .B2(_08741_),
    .Y(_08742_));
 sky130_vsdinv _25401_ (.A(_08514_),
    .Y(_08743_));
 sky130_fd_sc_hd__o21ai_4 _25402_ (.A1(_08455_),
    .A2(_08743_),
    .B1(_08456_),
    .Y(_08744_));
 sky130_fd_sc_hd__a21oi_2 _25403_ (.A1(_08740_),
    .A2(_08742_),
    .B1(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__nand3_4 _25404_ (.A(_08744_),
    .B(_08740_),
    .C(_08742_),
    .Y(_08746_));
 sky130_vsdinv _25405_ (.A(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__nor2_1 _25406_ (.A(_08484_),
    .B(_08505_),
    .Y(_08748_));
 sky130_fd_sc_hd__a21o_4 _25407_ (.A1(_08504_),
    .A2(_08486_),
    .B1(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__o21bai_4 _25408_ (.A1(_08458_),
    .A2(_08510_),
    .B1_N(_08511_),
    .Y(_08750_));
 sky130_fd_sc_hd__xor2_4 _25409_ (.A(_08749_),
    .B(_08750_),
    .X(_08751_));
 sky130_fd_sc_hd__o21bai_4 _25410_ (.A1(_08745_),
    .A2(_08747_),
    .B1_N(_08751_),
    .Y(_08752_));
 sky130_fd_sc_hd__a21o_1 _25411_ (.A1(_08740_),
    .A2(_08742_),
    .B1(_08744_),
    .X(_08753_));
 sky130_fd_sc_hd__nand3_4 _25412_ (.A(_08753_),
    .B(_08751_),
    .C(_08746_),
    .Y(_08754_));
 sky130_fd_sc_hd__or2b_1 _25413_ (.A(_08530_),
    .B_N(_08531_),
    .X(_08755_));
 sky130_fd_sc_hd__a21oi_2 _25414_ (.A1(_08515_),
    .A2(_08516_),
    .B1(_08520_),
    .Y(_08756_));
 sky130_fd_sc_hd__o21ai_4 _25415_ (.A1(_08755_),
    .A2(_08756_),
    .B1(_08521_),
    .Y(_08757_));
 sky130_fd_sc_hd__a21oi_2 _25416_ (.A1(_08752_),
    .A2(_08754_),
    .B1(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__nand3_4 _25417_ (.A(_08752_),
    .B(_08757_),
    .C(_08754_),
    .Y(_08759_));
 sky130_vsdinv _25418_ (.A(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__nand2_4 _25419_ (.A(_08531_),
    .B(_08524_),
    .Y(_08761_));
 sky130_fd_sc_hd__o21bai_4 _25420_ (.A1(_08758_),
    .A2(_08760_),
    .B1_N(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__a21o_2 _25421_ (.A1(_08752_),
    .A2(_08754_),
    .B1(_08757_),
    .X(_08763_));
 sky130_fd_sc_hd__nand3_4 _25422_ (.A(_08763_),
    .B(_08759_),
    .C(_08761_),
    .Y(_08764_));
 sky130_vsdinv _25423_ (.A(_08541_),
    .Y(_08765_));
 sky130_fd_sc_hd__a21oi_2 _25424_ (.A1(_08539_),
    .A2(_08534_),
    .B1(_08536_),
    .Y(_08766_));
 sky130_fd_sc_hd__o21ai_4 _25425_ (.A1(_08765_),
    .A2(_08766_),
    .B1(_08540_),
    .Y(_08767_));
 sky130_fd_sc_hd__a21oi_4 _25426_ (.A1(_08762_),
    .A2(_08764_),
    .B1(_08767_),
    .Y(_08768_));
 sky130_fd_sc_hd__nand3_4 _25427_ (.A(_08762_),
    .B(_08767_),
    .C(_08764_),
    .Y(_08769_));
 sky130_fd_sc_hd__or2b_4 _25428_ (.A(_08768_),
    .B_N(_08769_),
    .X(_08770_));
 sky130_fd_sc_hd__a21boi_1 _25429_ (.A1(_08567_),
    .A2(_08545_),
    .B1_N(_08546_),
    .Y(_08771_));
 sky130_fd_sc_hd__xor2_1 _25430_ (.A(_08770_),
    .B(_08771_),
    .X(_02652_));
 sky130_fd_sc_hd__a21boi_1 _25431_ (.A1(_08611_),
    .A2(_08586_),
    .B1_N(_08585_),
    .Y(_08772_));
 sky130_fd_sc_hd__nor2_1 _25432_ (.A(_08575_),
    .B(_08580_),
    .Y(_08773_));
 sky130_fd_sc_hd__o21ba_1 _25433_ (.A1(_08574_),
    .A2(_08581_),
    .B1_N(_08773_),
    .X(_08774_));
 sky130_fd_sc_hd__or2b_1 _25434_ (.A(_08713_),
    .B_N(_08704_),
    .X(_08775_));
 sky130_fd_sc_hd__o21ai_2 _25435_ (.A1(_08712_),
    .A2(_08705_),
    .B1(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__o21a_2 _25436_ (.A1(_08576_),
    .A2(_08579_),
    .B1(_08577_),
    .X(_08777_));
 sky130_fd_sc_hd__a2bb2oi_4 _25437_ (.A1_N(_14321_),
    .A2_N(_08700_),
    .B1(_08698_),
    .B2(_08702_),
    .Y(_08778_));
 sky130_fd_sc_hd__clkbuf_2 _25438_ (.A(\pcpi_mul.rs1[28] ),
    .X(_08779_));
 sky130_fd_sc_hd__and2_2 _25439_ (.A(_04998_),
    .B(_08779_),
    .X(_08780_));
 sky130_fd_sc_hd__nand3_4 _25440_ (.A(_05126_),
    .B(_05164_),
    .C(_07568_),
    .Y(_08781_));
 sky130_fd_sc_hd__clkbuf_4 _25441_ (.A(\pcpi_mul.rs1[27] ),
    .X(_08782_));
 sky130_fd_sc_hd__a22o_2 _25442_ (.A1(_05126_),
    .A2(_07476_),
    .B1(_05064_),
    .B2(_08782_),
    .X(_08783_));
 sky130_fd_sc_hd__o21ai_4 _25443_ (.A1(_14297_),
    .A2(_08781_),
    .B1(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__xor2_4 _25444_ (.A(_08780_),
    .B(_08784_),
    .X(_08785_));
 sky130_fd_sc_hd__xnor2_4 _25445_ (.A(_08778_),
    .B(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__xor2_4 _25446_ (.A(_08777_),
    .B(_08786_),
    .X(_08787_));
 sky130_fd_sc_hd__xnor2_1 _25447_ (.A(_08776_),
    .B(_08787_),
    .Y(_08788_));
 sky130_fd_sc_hd__xor2_1 _25448_ (.A(_08774_),
    .B(_08788_),
    .X(_08789_));
 sky130_vsdinv _25449_ (.A(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__and2_1 _25450_ (.A(_08582_),
    .B(_08573_),
    .X(_08791_));
 sky130_fd_sc_hd__o21ba_1 _25451_ (.A1(_08571_),
    .A2(_08583_),
    .B1_N(_08791_),
    .X(_08792_));
 sky130_fd_sc_hd__nor2_1 _25452_ (.A(_08790_),
    .B(_08792_),
    .Y(_08793_));
 sky130_vsdinv _25453_ (.A(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__nand2_2 _25454_ (.A(_08792_),
    .B(_08790_),
    .Y(_08795_));
 sky130_fd_sc_hd__nand3b_2 _25455_ (.A_N(_08599_),
    .B(_14084_),
    .C(_08482_),
    .Y(_08796_));
 sky130_fd_sc_hd__o31a_4 _25456_ (.A1(_14091_),
    .A2(_14277_),
    .A3(_08598_),
    .B1(_08796_),
    .X(_08797_));
 sky130_fd_sc_hd__nor2_1 _25457_ (.A(_08602_),
    .B(_08607_),
    .Y(_08798_));
 sky130_fd_sc_hd__o21bai_4 _25458_ (.A1(_08600_),
    .A2(_08608_),
    .B1_N(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__and2_2 _25459_ (.A(_14084_),
    .B(_08588_),
    .X(_08800_));
 sky130_fd_sc_hd__nand2_2 _25460_ (.A(_12776_),
    .B(\pcpi_mul.rs2[2] ),
    .Y(_08801_));
 sky130_fd_sc_hd__xnor2_4 _25461_ (.A(_08598_),
    .B(_08801_),
    .Y(_08802_));
 sky130_fd_sc_hd__xor2_4 _25462_ (.A(_08800_),
    .B(_08802_),
    .X(_08803_));
 sky130_fd_sc_hd__a21boi_4 _25463_ (.A1(_08601_),
    .A2(_08605_),
    .B1_N(_08603_),
    .Y(_08804_));
 sky130_fd_sc_hd__or4_4 _25464_ (.A(_14075_),
    .B(_14077_),
    .C(_14279_),
    .D(_14285_),
    .X(_08805_));
 sky130_fd_sc_hd__clkbuf_4 _25465_ (.A(_08078_),
    .X(_08806_));
 sky130_fd_sc_hd__a22o_2 _25466_ (.A1(_06159_),
    .A2(_08488_),
    .B1(_08604_),
    .B2(_08806_),
    .X(_08807_));
 sky130_fd_sc_hd__nand2_2 _25467_ (.A(_08805_),
    .B(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__xor2_4 _25468_ (.A(_08498_),
    .B(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__xnor2_4 _25469_ (.A(_08804_),
    .B(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__xor2_4 _25470_ (.A(_08803_),
    .B(_08810_),
    .X(_08811_));
 sky130_fd_sc_hd__xnor2_4 _25471_ (.A(_08799_),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__xor2_4 _25472_ (.A(_08797_),
    .B(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__a21o_1 _25473_ (.A1(_08794_),
    .A2(_08795_),
    .B1(_08813_),
    .X(_08814_));
 sky130_fd_sc_hd__nand3b_4 _25474_ (.A_N(_08793_),
    .B(_08813_),
    .C(_08795_),
    .Y(_08815_));
 sky130_fd_sc_hd__and2b_1 _25475_ (.A_N(_08697_),
    .B(_08731_),
    .X(_08816_));
 sky130_fd_sc_hd__o21bai_4 _25476_ (.A1(_08694_),
    .A2(_08732_),
    .B1_N(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__a21o_1 _25477_ (.A1(_08814_),
    .A2(_08815_),
    .B1(_08817_),
    .X(_08818_));
 sky130_fd_sc_hd__nand3_4 _25478_ (.A(_08814_),
    .B(_08817_),
    .C(_08815_),
    .Y(_08819_));
 sky130_fd_sc_hd__nand3b_4 _25479_ (.A_N(_08772_),
    .B(_08818_),
    .C(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__a21bo_2 _25480_ (.A1(_08818_),
    .A2(_08819_),
    .B1_N(_08772_),
    .X(_08821_));
 sky130_fd_sc_hd__o21a_2 _25481_ (.A1(_08625_),
    .A2(_08630_),
    .B1(_08626_),
    .X(_08822_));
 sky130_fd_sc_hd__a2bb2oi_4 _25482_ (.A1_N(_14429_),
    .A2_N(_08638_),
    .B1(_08635_),
    .B2(_08639_),
    .Y(_08823_));
 sky130_fd_sc_hd__nand2_4 _25483_ (.A(_08400_),
    .B(_05311_),
    .Y(_08824_));
 sky130_fd_sc_hd__or4_4 _25484_ (.A(_08402_),
    .B(_13990_),
    .C(_06127_),
    .D(_05998_),
    .X(_08825_));
 sky130_fd_sc_hd__a22o_1 _25485_ (.A1(_08404_),
    .A2(_05228_),
    .B1(_08405_),
    .B2(_05237_),
    .X(_08826_));
 sky130_fd_sc_hd__nand2_2 _25486_ (.A(_08825_),
    .B(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__xnor2_4 _25487_ (.A(_08824_),
    .B(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__xnor2_4 _25488_ (.A(_08823_),
    .B(_08828_),
    .Y(_08829_));
 sky130_fd_sc_hd__xor2_4 _25489_ (.A(_08822_),
    .B(_08829_),
    .X(_08830_));
 sky130_fd_sc_hd__or2b_1 _25490_ (.A(_08650_),
    .B_N(_08643_),
    .X(_08831_));
 sky130_fd_sc_hd__o21ai_2 _25491_ (.A1(_08641_),
    .A2(_08651_),
    .B1(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__and2_2 _25492_ (.A(_07358_),
    .B(_05819_),
    .X(_08833_));
 sky130_fd_sc_hd__nand3_4 _25493_ (.A(_08374_),
    .B(_08375_),
    .C(_05039_),
    .Y(_08834_));
 sky130_fd_sc_hd__a22o_2 _25494_ (.A1(_07961_),
    .A2(_05032_),
    .B1(_13977_),
    .B2(_05041_),
    .X(_08835_));
 sky130_fd_sc_hd__o21ai_4 _25495_ (.A1(_05057_),
    .A2(_08834_),
    .B1(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__xor2_4 _25496_ (.A(_08833_),
    .B(_08836_),
    .X(_08837_));
 sky130_fd_sc_hd__nand3b_2 _25497_ (.A_N(_08647_),
    .B(_08526_),
    .C(_14449_),
    .Y(_08838_));
 sky130_fd_sc_hd__o31ai_4 _25498_ (.A1(_13966_),
    .A2(_05178_),
    .A3(_08649_),
    .B1(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__and2_2 _25499_ (.A(_08644_),
    .B(_04927_),
    .X(_08840_));
 sky130_fd_sc_hd__nand2_2 _25500_ (.A(_08646_),
    .B(_05051_),
    .Y(_08841_));
 sky130_fd_sc_hd__and2b_1 _25501_ (.A_N(_04988_),
    .B(_08383_),
    .X(_08842_));
 sky130_fd_sc_hd__xor2_4 _25502_ (.A(_08841_),
    .B(_08842_),
    .X(_08843_));
 sky130_fd_sc_hd__xor2_4 _25503_ (.A(_08840_),
    .B(_08843_),
    .X(_08844_));
 sky130_fd_sc_hd__xor2_4 _25504_ (.A(_08839_),
    .B(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__xor2_4 _25505_ (.A(_08837_),
    .B(_08845_),
    .X(_08846_));
 sky130_fd_sc_hd__xnor2_2 _25506_ (.A(_08832_),
    .B(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__xnor2_2 _25507_ (.A(_08830_),
    .B(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__nand2_2 _25508_ (.A(_08653_),
    .B(_08652_),
    .Y(_08849_));
 sky130_fd_sc_hd__or2b_2 _25509_ (.A(_08654_),
    .B_N(_08633_),
    .X(_08850_));
 sky130_fd_sc_hd__nand3b_4 _25510_ (.A_N(_08848_),
    .B(_08849_),
    .C(_08850_),
    .Y(_08851_));
 sky130_fd_sc_hd__nand2_1 _25511_ (.A(_08850_),
    .B(_08849_),
    .Y(_08852_));
 sky130_fd_sc_hd__nand2_4 _25512_ (.A(_08852_),
    .B(_08848_),
    .Y(_08853_));
 sky130_fd_sc_hd__nor2_1 _25513_ (.A(_08666_),
    .B(_08675_),
    .Y(_08854_));
 sky130_fd_sc_hd__o21ba_2 _25514_ (.A1(_08665_),
    .A2(_08676_),
    .B1_N(_08854_),
    .X(_08855_));
 sky130_fd_sc_hd__and2_2 _25515_ (.A(_06060_),
    .B(_05778_),
    .X(_08856_));
 sky130_fd_sc_hd__buf_6 _25516_ (.A(_08662_),
    .X(_08857_));
 sky130_fd_sc_hd__nand3_4 _25517_ (.A(_08857_),
    .B(_08423_),
    .C(_05692_),
    .Y(_08858_));
 sky130_fd_sc_hd__buf_6 _25518_ (.A(_14015_),
    .X(_08859_));
 sky130_fd_sc_hd__a22o_2 _25519_ (.A1(_08660_),
    .A2(_05611_),
    .B1(_08859_),
    .B2(_05700_),
    .X(_08860_));
 sky130_fd_sc_hd__o21ai_4 _25520_ (.A1(_14374_),
    .A2(_08858_),
    .B1(_08860_),
    .Y(_08861_));
 sky130_fd_sc_hd__xor2_4 _25521_ (.A(_08856_),
    .B(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__o21a_2 _25522_ (.A1(_14395_),
    .A2(_08670_),
    .B1(_08674_),
    .X(_08863_));
 sky130_fd_sc_hd__buf_4 _25523_ (.A(_07979_),
    .X(_08864_));
 sky130_fd_sc_hd__a22o_1 _25524_ (.A1(_08431_),
    .A2(_05497_),
    .B1(_08864_),
    .B2(_08264_),
    .X(_08865_));
 sky130_fd_sc_hd__nand3_4 _25525_ (.A(_08431_),
    .B(_08432_),
    .C(_05413_),
    .Y(_08866_));
 sky130_fd_sc_hd__or2b_1 _25526_ (.A(_08866_),
    .B_N(_05505_),
    .X(_08867_));
 sky130_fd_sc_hd__o2bb2ai_1 _25527_ (.A1_N(_08865_),
    .A2_N(_08867_),
    .B1(_14006_),
    .B2(_06409_),
    .Y(_08868_));
 sky130_fd_sc_hd__o2111ai_4 _25528_ (.A1(_14389_),
    .A2(_08866_),
    .B1(_06471_),
    .C1(_06161_),
    .D1(_08865_),
    .Y(_08869_));
 sky130_fd_sc_hd__nand2_4 _25529_ (.A(_08868_),
    .B(_08869_),
    .Y(_08870_));
 sky130_fd_sc_hd__xnor2_4 _25530_ (.A(_08863_),
    .B(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__xor2_4 _25531_ (.A(_08862_),
    .B(_08871_),
    .X(_08872_));
 sky130_fd_sc_hd__nor2_1 _25532_ (.A(_08624_),
    .B(_08631_),
    .Y(_08873_));
 sky130_fd_sc_hd__o21bai_4 _25533_ (.A1(_08623_),
    .A2(_08632_),
    .B1_N(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__xnor2_4 _25534_ (.A(_08872_),
    .B(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__xor2_4 _25535_ (.A(_08855_),
    .B(_08875_),
    .X(_08876_));
 sky130_fd_sc_hd__a21oi_1 _25536_ (.A1(_08851_),
    .A2(_08853_),
    .B1(_08876_),
    .Y(_08877_));
 sky130_vsdinv _25537_ (.A(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__nand3_4 _25538_ (.A(_08851_),
    .B(_08876_),
    .C(_08853_),
    .Y(_08879_));
 sky130_fd_sc_hd__o21ai_4 _25539_ (.A1(_08656_),
    .A2(_08682_),
    .B1(_08683_),
    .Y(_08880_));
 sky130_fd_sc_hd__a21oi_4 _25540_ (.A1(_08878_),
    .A2(_08879_),
    .B1(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__o211a_1 _25541_ (.A1(_08685_),
    .A2(_08684_),
    .B1(_08879_),
    .C1(_08878_),
    .X(_08882_));
 sky130_fd_sc_hd__nand2_1 _25542_ (.A(_08729_),
    .B(_08717_),
    .Y(_08883_));
 sky130_fd_sc_hd__o21a_2 _25543_ (.A1(_08715_),
    .A2(_08730_),
    .B1(_08883_),
    .X(_08884_));
 sky130_fd_sc_hd__buf_2 _25544_ (.A(_07044_),
    .X(_08885_));
 sky130_fd_sc_hd__and2_2 _25545_ (.A(_05206_),
    .B(_08885_),
    .X(_08886_));
 sky130_fd_sc_hd__nand3_4 _25546_ (.A(_08333_),
    .B(_05274_),
    .C(_08330_),
    .Y(_08887_));
 sky130_fd_sc_hd__a22o_2 _25547_ (.A1(_08333_),
    .A2(_07206_),
    .B1(_05364_),
    .B2(_08085_),
    .X(_08888_));
 sky130_fd_sc_hd__o21ai_4 _25548_ (.A1(_14315_),
    .A2(_08887_),
    .B1(_08888_),
    .Y(_08889_));
 sky130_fd_sc_hd__xnor2_4 _25549_ (.A(_08886_),
    .B(_08889_),
    .Y(_08890_));
 sky130_fd_sc_hd__o21a_4 _25550_ (.A1(_14340_),
    .A2(_08707_),
    .B1(_08711_),
    .X(_08891_));
 sky130_fd_sc_hd__a22o_1 _25551_ (.A1(_07655_),
    .A2(_06296_),
    .B1(_05531_),
    .B2(_07048_),
    .X(_08892_));
 sky130_fd_sc_hd__nand3_4 _25552_ (.A(_07655_),
    .B(_05531_),
    .C(_07046_),
    .Y(_08893_));
 sky130_fd_sc_hd__or2b_1 _25553_ (.A(_08893_),
    .B_N(_06450_),
    .X(_08894_));
 sky130_fd_sc_hd__o2bb2ai_1 _25554_ (.A1_N(_08892_),
    .A2_N(_08894_),
    .B1(_14048_),
    .B2(_14327_),
    .Y(_08895_));
 sky130_fd_sc_hd__o2111ai_4 _25555_ (.A1(_14333_),
    .A2(_08893_),
    .B1(_08710_),
    .C1(_06940_),
    .D1(_08892_),
    .Y(_08896_));
 sky130_fd_sc_hd__nand2_4 _25556_ (.A(_08895_),
    .B(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__xnor2_4 _25557_ (.A(_08891_),
    .B(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__xnor2_4 _25558_ (.A(_08890_),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__nor2_1 _25559_ (.A(_08719_),
    .B(_08727_),
    .Y(_08900_));
 sky130_fd_sc_hd__o21bai_4 _25560_ (.A1(_08718_),
    .A2(_08728_),
    .B1_N(_08900_),
    .Y(_08901_));
 sky130_fd_sc_hd__o21a_4 _25561_ (.A1(_14361_),
    .A2(_08723_),
    .B1(_08726_),
    .X(_08902_));
 sky130_fd_sc_hd__a2bb2oi_4 _25562_ (.A1_N(_08210_),
    .A2_N(_08661_),
    .B1(_08659_),
    .B2(_08663_),
    .Y(_08903_));
 sky130_fd_sc_hd__a22o_1 _25563_ (.A1(_05943_),
    .A2(_06029_),
    .B1(_05944_),
    .B2(_06037_),
    .X(_08904_));
 sky130_fd_sc_hd__nand3_4 _25564_ (.A(_06349_),
    .B(_08357_),
    .C(_05912_),
    .Y(_08905_));
 sky130_fd_sc_hd__or2b_1 _25565_ (.A(_08905_),
    .B_N(_06155_),
    .X(_08906_));
 sky130_fd_sc_hd__o2bb2ai_1 _25566_ (.A1_N(_08904_),
    .A2_N(_08906_),
    .B1(_14032_),
    .B2(_06293_),
    .Y(_08907_));
 sky130_fd_sc_hd__o2111ai_4 _25567_ (.A1(_14353_),
    .A2(_08905_),
    .B1(_05939_),
    .C1(_08342_),
    .D1(_08904_),
    .Y(_08908_));
 sky130_fd_sc_hd__nand2_4 _25568_ (.A(_08907_),
    .B(_08908_),
    .Y(_08909_));
 sky130_fd_sc_hd__xnor2_4 _25569_ (.A(_08903_),
    .B(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__xor2_4 _25570_ (.A(_08902_),
    .B(_08910_),
    .X(_08911_));
 sky130_fd_sc_hd__xnor2_4 _25571_ (.A(_08901_),
    .B(_08911_),
    .Y(_08912_));
 sky130_fd_sc_hd__xnor2_4 _25572_ (.A(_08899_),
    .B(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__and2_1 _25573_ (.A(_08679_),
    .B(_08677_),
    .X(_08914_));
 sky130_fd_sc_hd__o21ba_2 _25574_ (.A1(_08658_),
    .A2(_08680_),
    .B1_N(_08914_),
    .X(_08915_));
 sky130_fd_sc_hd__xor2_4 _25575_ (.A(_08913_),
    .B(_08915_),
    .X(_08916_));
 sky130_fd_sc_hd__xor2_4 _25576_ (.A(_08884_),
    .B(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__o21bai_4 _25577_ (.A1(_08881_),
    .A2(_08882_),
    .B1_N(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__nand3b_4 _25578_ (.A_N(_08877_),
    .B(_08879_),
    .C(_08880_),
    .Y(_08919_));
 sky130_fd_sc_hd__nand3b_4 _25579_ (.A_N(_08881_),
    .B(_08917_),
    .C(_08919_),
    .Y(_08920_));
 sky130_vsdinv _25580_ (.A(_08733_),
    .Y(_08921_));
 sky130_fd_sc_hd__o21bai_4 _25581_ (.A1(_08921_),
    .A2(_08688_),
    .B1_N(_08690_),
    .Y(_08922_));
 sky130_fd_sc_hd__a21o_1 _25582_ (.A1(_08918_),
    .A2(_08920_),
    .B1(_08922_),
    .X(_08923_));
 sky130_fd_sc_hd__nand3_4 _25583_ (.A(_08918_),
    .B(_08920_),
    .C(_08922_),
    .Y(_08924_));
 sky130_fd_sc_hd__a22oi_4 _25584_ (.A1(_08820_),
    .A2(_08821_),
    .B1(_08923_),
    .B2(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__a21oi_4 _25585_ (.A1(_08918_),
    .A2(_08920_),
    .B1(_08922_),
    .Y(_08926_));
 sky130_fd_sc_hd__nand2_2 _25586_ (.A(_08821_),
    .B(_08820_),
    .Y(_08927_));
 sky130_fd_sc_hd__nor3b_4 _25587_ (.A(_08926_),
    .B(_08927_),
    .C_N(_08924_),
    .Y(_08928_));
 sky130_fd_sc_hd__o31ai_4 _25588_ (.A1(_08619_),
    .A2(_08620_),
    .A3(_08737_),
    .B1(_08739_),
    .Y(_08929_));
 sky130_fd_sc_hd__o21bai_4 _25589_ (.A1(_08925_),
    .A2(_08928_),
    .B1_N(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__a22o_1 _25590_ (.A1(_08820_),
    .A2(_08821_),
    .B1(_08923_),
    .B2(_08924_),
    .X(_08931_));
 sky130_fd_sc_hd__nand3b_2 _25591_ (.A_N(_08927_),
    .B(_08924_),
    .C(_08923_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand3_4 _25592_ (.A(_08931_),
    .B(_08929_),
    .C(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__nor2_1 _25593_ (.A(_08591_),
    .B(_08610_),
    .Y(_08934_));
 sky130_fd_sc_hd__a21o_4 _25594_ (.A1(_08609_),
    .A2(_08593_),
    .B1(_08934_),
    .X(_08935_));
 sky130_fd_sc_hd__nand3b_4 _25595_ (.A_N(_08618_),
    .B(_08616_),
    .C(_08617_),
    .Y(_08936_));
 sky130_fd_sc_hd__nand2_2 _25596_ (.A(_08936_),
    .B(_08617_),
    .Y(_08937_));
 sky130_fd_sc_hd__xor2_4 _25597_ (.A(_08935_),
    .B(_08937_),
    .X(_08938_));
 sky130_fd_sc_hd__a21oi_4 _25598_ (.A1(_08930_),
    .A2(_08933_),
    .B1(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__nand3_4 _25599_ (.A(_08930_),
    .B(_08938_),
    .C(_08933_),
    .Y(_08940_));
 sky130_vsdinv _25600_ (.A(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__a21o_1 _25601_ (.A1(_08753_),
    .A2(_08751_),
    .B1(_08747_),
    .X(_08942_));
 sky130_fd_sc_hd__o21bai_4 _25602_ (.A1(_08939_),
    .A2(_08941_),
    .B1_N(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__a21o_1 _25603_ (.A1(_08930_),
    .A2(_08933_),
    .B1(_08938_),
    .X(_08944_));
 sky130_fd_sc_hd__nand3_4 _25604_ (.A(_08944_),
    .B(_08942_),
    .C(_08940_),
    .Y(_08945_));
 sky130_fd_sc_hd__and2_2 _25605_ (.A(_08750_),
    .B(_08749_),
    .X(_08946_));
 sky130_fd_sc_hd__a21oi_4 _25606_ (.A1(_08943_),
    .A2(_08945_),
    .B1(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__nand3_4 _25607_ (.A(_08943_),
    .B(_08946_),
    .C(_08945_),
    .Y(_08948_));
 sky130_vsdinv _25608_ (.A(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__a21oi_4 _25609_ (.A1(_08763_),
    .A2(_08761_),
    .B1(_08760_),
    .Y(_08950_));
 sky130_fd_sc_hd__o21ai_1 _25610_ (.A1(_08947_),
    .A2(_08949_),
    .B1(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__a21o_1 _25611_ (.A1(_08763_),
    .A2(_08761_),
    .B1(_08760_),
    .X(_08952_));
 sky130_fd_sc_hd__nand2_1 _25612_ (.A(_08943_),
    .B(_08945_),
    .Y(_08953_));
 sky130_vsdinv _25613_ (.A(_08946_),
    .Y(_08954_));
 sky130_fd_sc_hd__nand2_2 _25614_ (.A(_08953_),
    .B(_08954_),
    .Y(_08955_));
 sky130_fd_sc_hd__nand3_4 _25615_ (.A(_08952_),
    .B(_08955_),
    .C(_08948_),
    .Y(_08956_));
 sky130_fd_sc_hd__nand2_2 _25616_ (.A(_08951_),
    .B(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__nor2_8 _25617_ (.A(_08547_),
    .B(_08770_),
    .Y(_08958_));
 sky130_fd_sc_hd__a21oi_4 _25618_ (.A1(_08546_),
    .A2(_08769_),
    .B1(_08768_),
    .Y(_08959_));
 sky130_fd_sc_hd__a21oi_2 _25619_ (.A1(_08567_),
    .A2(_08958_),
    .B1(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__xor2_1 _25620_ (.A(_08957_),
    .B(_08960_),
    .X(_02653_));
 sky130_fd_sc_hd__nor2_1 _25621_ (.A(_08777_),
    .B(_08786_),
    .Y(_08961_));
 sky130_fd_sc_hd__o21ba_2 _25622_ (.A1(_08778_),
    .A2(_08785_),
    .B1_N(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__or2b_1 _25623_ (.A(_08898_),
    .B_N(_08890_),
    .X(_08963_));
 sky130_fd_sc_hd__o21ai_4 _25624_ (.A1(_08897_),
    .A2(_08891_),
    .B1(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__a2bb2oi_4 _25625_ (.A1_N(_14300_),
    .A2_N(_08781_),
    .B1(_08780_),
    .B2(_08783_),
    .Y(_08965_));
 sky130_fd_sc_hd__a2bb2oi_4 _25626_ (.A1_N(_08464_),
    .A2_N(_08887_),
    .B1(_08886_),
    .B2(_08888_),
    .Y(_08966_));
 sky130_fd_sc_hd__nand2_4 _25627_ (.A(_04998_),
    .B(_08488_),
    .Y(_08967_));
 sky130_fd_sc_hd__or4_4 _25628_ (.A(_14063_),
    .B(_14067_),
    .C(_14290_),
    .D(_14296_),
    .X(_08968_));
 sky130_fd_sc_hd__a22o_1 _25629_ (.A1(_05132_),
    .A2(_07485_),
    .B1(_05164_),
    .B2(_08779_),
    .X(_08969_));
 sky130_fd_sc_hd__nand2_2 _25630_ (.A(_08968_),
    .B(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__xnor2_4 _25631_ (.A(_08967_),
    .B(_08970_),
    .Y(_08971_));
 sky130_fd_sc_hd__xnor2_4 _25632_ (.A(_08966_),
    .B(_08971_),
    .Y(_08972_));
 sky130_fd_sc_hd__xor2_4 _25633_ (.A(_08965_),
    .B(_08972_),
    .X(_08973_));
 sky130_fd_sc_hd__xnor2_4 _25634_ (.A(_08964_),
    .B(_08973_),
    .Y(_08974_));
 sky130_fd_sc_hd__xor2_4 _25635_ (.A(_08962_),
    .B(_08974_),
    .X(_08975_));
 sky130_fd_sc_hd__and2_1 _25636_ (.A(_08787_),
    .B(_08776_),
    .X(_08976_));
 sky130_fd_sc_hd__o21ba_1 _25637_ (.A1(_08774_),
    .A2(_08788_),
    .B1_N(_08976_),
    .X(_08977_));
 sky130_fd_sc_hd__or2b_2 _25638_ (.A(_08975_),
    .B_N(_08977_),
    .X(_08978_));
 sky130_vsdinv _25639_ (.A(_08977_),
    .Y(_08979_));
 sky130_fd_sc_hd__nand2_2 _25640_ (.A(_08975_),
    .B(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__nand3_4 _25641_ (.A(_12781_),
    .B(_04886_),
    .C(_04878_),
    .Y(_08981_));
 sky130_fd_sc_hd__o31a_4 _25642_ (.A1(_14088_),
    .A2(_14277_),
    .A3(_08802_),
    .B1(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__nor2_1 _25643_ (.A(_08804_),
    .B(_08809_),
    .Y(_08983_));
 sky130_fd_sc_hd__o21bai_4 _25644_ (.A1(_08803_),
    .A2(_08810_),
    .B1_N(_08983_),
    .Y(_08984_));
 sky130_fd_sc_hd__nand2_4 _25645_ (.A(_12777_),
    .B(\pcpi_mul.rs2[3] ),
    .Y(_08985_));
 sky130_fd_sc_hd__xor2_4 _25646_ (.A(_08985_),
    .B(_08802_),
    .X(_08986_));
 sky130_fd_sc_hd__clkinv_4 _25647_ (.A(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__a21boi_4 _25648_ (.A1(_08601_),
    .A2(_08807_),
    .B1_N(_08805_),
    .Y(_08988_));
 sky130_fd_sc_hd__or4_4 _25649_ (.A(_14075_),
    .B(_14077_),
    .C(_14275_),
    .D(_14279_),
    .X(_08989_));
 sky130_fd_sc_hd__a22o_2 _25650_ (.A1(_05420_),
    .A2(_08480_),
    .B1(_08604_),
    .B2(_08492_),
    .X(_08990_));
 sky130_fd_sc_hd__nand2_4 _25651_ (.A(_08989_),
    .B(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__xor2_4 _25652_ (.A(_08601_),
    .B(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__xnor2_4 _25653_ (.A(_08988_),
    .B(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__xor2_4 _25654_ (.A(_08987_),
    .B(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__xnor2_4 _25655_ (.A(_08984_),
    .B(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__xor2_4 _25656_ (.A(_08982_),
    .B(_08995_),
    .X(_08996_));
 sky130_fd_sc_hd__a21o_1 _25657_ (.A1(_08978_),
    .A2(_08980_),
    .B1(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__nand3_4 _25658_ (.A(_08978_),
    .B(_08996_),
    .C(_08980_),
    .Y(_08998_));
 sky130_fd_sc_hd__and2b_1 _25659_ (.A_N(_08915_),
    .B(_08913_),
    .X(_08999_));
 sky130_fd_sc_hd__o21bai_4 _25660_ (.A1(_08884_),
    .A2(_08916_),
    .B1_N(_08999_),
    .Y(_09000_));
 sky130_fd_sc_hd__a21o_1 _25661_ (.A1(_08997_),
    .A2(_08998_),
    .B1(_09000_),
    .X(_09001_));
 sky130_fd_sc_hd__a21oi_1 _25662_ (.A1(_08795_),
    .A2(_08813_),
    .B1(_08793_),
    .Y(_09002_));
 sky130_vsdinv _25663_ (.A(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__nand3_4 _25664_ (.A(_08997_),
    .B(_09000_),
    .C(_08998_),
    .Y(_09004_));
 sky130_fd_sc_hd__nand3_4 _25665_ (.A(_09001_),
    .B(_09003_),
    .C(_09004_),
    .Y(_09005_));
 sky130_fd_sc_hd__a21o_2 _25666_ (.A1(_09001_),
    .A2(_09004_),
    .B1(_09003_),
    .X(_09006_));
 sky130_fd_sc_hd__nand2_2 _25667_ (.A(_08846_),
    .B(_08832_),
    .Y(_09007_));
 sky130_fd_sc_hd__or2b_2 _25668_ (.A(_08847_),
    .B_N(_08830_),
    .X(_09008_));
 sky130_fd_sc_hd__o21a_2 _25669_ (.A1(_08824_),
    .A2(_08827_),
    .B1(_08825_),
    .X(_09009_));
 sky130_fd_sc_hd__a2bb2oi_4 _25670_ (.A1_N(_14423_),
    .A2_N(_08834_),
    .B1(_08833_),
    .B2(_08835_),
    .Y(_09010_));
 sky130_fd_sc_hd__nand2_2 _25671_ (.A(_07106_),
    .B(_05414_),
    .Y(_09011_));
 sky130_fd_sc_hd__or4_4 _25672_ (.A(_08402_),
    .B(_13989_),
    .C(_14399_),
    .D(_14404_),
    .X(_09012_));
 sky130_fd_sc_hd__a22o_1 _25673_ (.A1(_07262_),
    .A2(_05516_),
    .B1(_07102_),
    .B2(_05614_),
    .X(_09013_));
 sky130_fd_sc_hd__nand2_2 _25674_ (.A(_09012_),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__xnor2_4 _25675_ (.A(_09011_),
    .B(_09014_),
    .Y(_09015_));
 sky130_fd_sc_hd__xnor2_4 _25676_ (.A(_09010_),
    .B(_09015_),
    .Y(_09016_));
 sky130_fd_sc_hd__xor2_2 _25677_ (.A(_09009_),
    .B(_09016_),
    .X(_09017_));
 sky130_fd_sc_hd__or2b_1 _25678_ (.A(_08844_),
    .B_N(_08839_),
    .X(_09018_));
 sky130_fd_sc_hd__o21ai_1 _25679_ (.A1(_08837_),
    .A2(_08845_),
    .B1(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__and2_2 _25680_ (.A(_07358_),
    .B(_05875_),
    .X(_09020_));
 sky130_fd_sc_hd__nand3_4 _25681_ (.A(_07961_),
    .B(_08375_),
    .C(_05041_),
    .Y(_09021_));
 sky130_fd_sc_hd__a22o_2 _25682_ (.A1(_13971_),
    .A2(_05099_),
    .B1(_13977_),
    .B2(_05101_),
    .X(_09022_));
 sky130_fd_sc_hd__o21ai_4 _25683_ (.A1(_05115_),
    .A2(_09021_),
    .B1(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__xor2_4 _25684_ (.A(_09020_),
    .B(_09023_),
    .X(_09024_));
 sky130_fd_sc_hd__buf_4 _25685_ (.A(_12804_),
    .X(_09025_));
 sky130_fd_sc_hd__nand3b_2 _25686_ (.A_N(_08841_),
    .B(_09025_),
    .C(_14443_),
    .Y(_09026_));
 sky130_fd_sc_hd__o31ai_4 _25687_ (.A1(_13966_),
    .A2(_05580_),
    .A3(_08843_),
    .B1(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__and2_2 _25688_ (.A(\pcpi_mul.rs2[30] ),
    .B(_05959_),
    .X(_09028_));
 sky130_fd_sc_hd__nand2_2 _25689_ (.A(_08646_),
    .B(_05111_),
    .Y(_09029_));
 sky130_fd_sc_hd__and2b_2 _25690_ (.A_N(_04948_),
    .B(\pcpi_mul.rs2[32] ),
    .X(_09030_));
 sky130_fd_sc_hd__xor2_4 _25691_ (.A(_09029_),
    .B(_09030_),
    .X(_09031_));
 sky130_fd_sc_hd__xor2_4 _25692_ (.A(_09028_),
    .B(_09031_),
    .X(_09032_));
 sky130_fd_sc_hd__xor2_4 _25693_ (.A(_09027_),
    .B(_09032_),
    .X(_09033_));
 sky130_fd_sc_hd__xor2_2 _25694_ (.A(_09024_),
    .B(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__xnor2_1 _25695_ (.A(_09019_),
    .B(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__xnor2_1 _25696_ (.A(_09017_),
    .B(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__a21bo_2 _25697_ (.A1(_09007_),
    .A2(_09008_),
    .B1_N(_09036_),
    .X(_09037_));
 sky130_fd_sc_hd__nand3b_4 _25698_ (.A_N(_09036_),
    .B(_09007_),
    .C(_09008_),
    .Y(_09038_));
 sky130_fd_sc_hd__nor2_1 _25699_ (.A(_08863_),
    .B(_08870_),
    .Y(_09039_));
 sky130_fd_sc_hd__o21ba_2 _25700_ (.A1(_08862_),
    .A2(_08871_),
    .B1_N(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__and2_2 _25701_ (.A(_06346_),
    .B(_06285_),
    .X(_09041_));
 sky130_fd_sc_hd__nand3_4 _25702_ (.A(_08422_),
    .B(_08859_),
    .C(_05770_),
    .Y(_09042_));
 sky130_fd_sc_hd__a22o_2 _25703_ (.A1(_08425_),
    .A2(_05700_),
    .B1(_08426_),
    .B2(_05778_),
    .X(_09043_));
 sky130_fd_sc_hd__o21ai_4 _25704_ (.A1(_14367_),
    .A2(_09042_),
    .B1(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__xor2_4 _25705_ (.A(_09041_),
    .B(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__o21a_2 _25706_ (.A1(_14390_),
    .A2(_08866_),
    .B1(_08869_),
    .X(_09046_));
 sky130_fd_sc_hd__a22o_1 _25707_ (.A1(_08667_),
    .A2(_08264_),
    .B1(_08864_),
    .B2(_06160_),
    .X(_09047_));
 sky130_fd_sc_hd__nand3_4 _25708_ (.A(_08269_),
    .B(_06647_),
    .C(_08264_),
    .Y(_09048_));
 sky130_fd_sc_hd__or2b_1 _25709_ (.A(_09048_),
    .B_N(_05513_),
    .X(_09049_));
 sky130_fd_sc_hd__o2bb2ai_1 _25710_ (.A1_N(_09047_),
    .A2_N(_09049_),
    .B1(_07123_),
    .B2(_08210_),
    .Y(_09050_));
 sky130_fd_sc_hd__o2111ai_4 _25711_ (.A1(_14384_),
    .A2(_09048_),
    .B1(_06471_),
    .C1(_05611_),
    .D1(_09047_),
    .Y(_09051_));
 sky130_fd_sc_hd__nand2_4 _25712_ (.A(_09050_),
    .B(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__xnor2_4 _25713_ (.A(_09046_),
    .B(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__xor2_4 _25714_ (.A(_09045_),
    .B(_09053_),
    .X(_09054_));
 sky130_fd_sc_hd__nor2_1 _25715_ (.A(_08823_),
    .B(_08828_),
    .Y(_09055_));
 sky130_fd_sc_hd__o21bai_4 _25716_ (.A1(_08822_),
    .A2(_08829_),
    .B1_N(_09055_),
    .Y(_09056_));
 sky130_fd_sc_hd__xnor2_4 _25717_ (.A(_09054_),
    .B(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__xor2_4 _25718_ (.A(_09040_),
    .B(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__a21oi_2 _25719_ (.A1(_09037_),
    .A2(_09038_),
    .B1(_09058_),
    .Y(_09059_));
 sky130_vsdinv _25720_ (.A(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__nand3_4 _25721_ (.A(_09037_),
    .B(_09058_),
    .C(_09038_),
    .Y(_09061_));
 sky130_fd_sc_hd__nand2_4 _25722_ (.A(_08879_),
    .B(_08853_),
    .Y(_09062_));
 sky130_fd_sc_hd__a21o_1 _25723_ (.A1(_09060_),
    .A2(_09061_),
    .B1(_09062_),
    .X(_09063_));
 sky130_fd_sc_hd__nand3b_4 _25724_ (.A_N(_09059_),
    .B(_09061_),
    .C(_09062_),
    .Y(_09064_));
 sky130_fd_sc_hd__and2_2 _25725_ (.A(_05206_),
    .B(_07569_),
    .X(_09065_));
 sky130_fd_sc_hd__nand3_4 _25726_ (.A(_05362_),
    .B(_05364_),
    .C(_08085_),
    .Y(_09066_));
 sky130_fd_sc_hd__a22o_2 _25727_ (.A1(_05362_),
    .A2(_07198_),
    .B1(_05364_),
    .B2(_07467_),
    .X(_09067_));
 sky130_fd_sc_hd__o21ai_4 _25728_ (.A1(_14309_),
    .A2(_09066_),
    .B1(_09067_),
    .Y(_09068_));
 sky130_fd_sc_hd__xnor2_4 _25729_ (.A(_09065_),
    .B(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__o21a_4 _25730_ (.A1(_07214_),
    .A2(_08893_),
    .B1(_08896_),
    .X(_09070_));
 sky130_fd_sc_hd__clkbuf_4 _25731_ (.A(_05637_),
    .X(_09071_));
 sky130_fd_sc_hd__a22o_1 _25732_ (.A1(_07281_),
    .A2(_07048_),
    .B1(_09071_),
    .B2(_06596_),
    .X(_09072_));
 sky130_fd_sc_hd__nand3_4 _25733_ (.A(_05955_),
    .B(_08199_),
    .C(_14331_),
    .Y(_09073_));
 sky130_fd_sc_hd__or2b_1 _25734_ (.A(_09073_),
    .B_N(_07033_),
    .X(_09074_));
 sky130_fd_sc_hd__o2bb2ai_1 _25735_ (.A1_N(_09072_),
    .A2_N(_09074_),
    .B1(_14047_),
    .B2(_08699_),
    .Y(_09075_));
 sky130_fd_sc_hd__o2111ai_4 _25736_ (.A1(_14326_),
    .A2(_09073_),
    .B1(_08710_),
    .C1(_07206_),
    .D1(_09072_),
    .Y(_09076_));
 sky130_fd_sc_hd__nand2_4 _25737_ (.A(_09075_),
    .B(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__xnor2_4 _25738_ (.A(_09070_),
    .B(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__xnor2_4 _25739_ (.A(_09069_),
    .B(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__nor2_1 _25740_ (.A(_08903_),
    .B(_08909_),
    .Y(_09080_));
 sky130_fd_sc_hd__o21bai_4 _25741_ (.A1(_08902_),
    .A2(_08910_),
    .B1_N(_09080_),
    .Y(_09081_));
 sky130_fd_sc_hd__o21a_4 _25742_ (.A1(_14354_),
    .A2(_08905_),
    .B1(_08908_),
    .X(_09082_));
 sky130_fd_sc_hd__a2bb2oi_4 _25743_ (.A1_N(_14373_),
    .A2_N(_08858_),
    .B1(_08856_),
    .B2(_08860_),
    .Y(_09083_));
 sky130_fd_sc_hd__nand2_4 _25744_ (.A(_05939_),
    .B(_07747_),
    .Y(_09084_));
 sky130_fd_sc_hd__or4_4 _25745_ (.A(_14024_),
    .B(_14028_),
    .C(_14345_),
    .D(_14351_),
    .X(_09085_));
 sky130_fd_sc_hd__a22o_1 _25746_ (.A1(_05941_),
    .A2(_06037_),
    .B1(_05944_),
    .B2(_06165_),
    .X(_09086_));
 sky130_fd_sc_hd__nand2_2 _25747_ (.A(_09085_),
    .B(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__xnor2_4 _25748_ (.A(_09084_),
    .B(_09087_),
    .Y(_09088_));
 sky130_fd_sc_hd__xnor2_4 _25749_ (.A(_09083_),
    .B(_09088_),
    .Y(_09089_));
 sky130_fd_sc_hd__xor2_4 _25750_ (.A(_09082_),
    .B(_09089_),
    .X(_09090_));
 sky130_fd_sc_hd__xnor2_1 _25751_ (.A(_09081_),
    .B(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__xnor2_1 _25752_ (.A(_09079_),
    .B(_09091_),
    .Y(_09092_));
 sky130_fd_sc_hd__and2_1 _25753_ (.A(_08874_),
    .B(_08872_),
    .X(_09093_));
 sky130_fd_sc_hd__o21ba_1 _25754_ (.A1(_08855_),
    .A2(_08875_),
    .B1_N(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__or2b_2 _25755_ (.A(_09092_),
    .B_N(_09094_),
    .X(_09095_));
 sky130_fd_sc_hd__or2b_2 _25756_ (.A(_09094_),
    .B_N(_09092_),
    .X(_09096_));
 sky130_fd_sc_hd__or2b_1 _25757_ (.A(_08912_),
    .B_N(_08899_),
    .X(_09097_));
 sky130_fd_sc_hd__a21boi_1 _25758_ (.A1(_08911_),
    .A2(_08901_),
    .B1_N(_09097_),
    .Y(_09098_));
 sky130_vsdinv _25759_ (.A(_09098_),
    .Y(_09099_));
 sky130_fd_sc_hd__a21o_1 _25760_ (.A1(_09095_),
    .A2(_09096_),
    .B1(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__nand3_4 _25761_ (.A(_09095_),
    .B(_09096_),
    .C(_09099_),
    .Y(_09101_));
 sky130_fd_sc_hd__nand2_4 _25762_ (.A(_09100_),
    .B(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__a21boi_2 _25763_ (.A1(_09063_),
    .A2(_09064_),
    .B1_N(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__a21oi_4 _25764_ (.A1(_09060_),
    .A2(_09061_),
    .B1(_09062_),
    .Y(_09104_));
 sky130_fd_sc_hd__nor3b_4 _25765_ (.A(_09102_),
    .B(_09104_),
    .C_N(_09064_),
    .Y(_09105_));
 sky130_vsdinv _25766_ (.A(_08917_),
    .Y(_09106_));
 sky130_fd_sc_hd__o21ai_4 _25767_ (.A1(_08881_),
    .A2(_09106_),
    .B1(_08919_),
    .Y(_09107_));
 sky130_fd_sc_hd__o21bai_4 _25768_ (.A1(_09103_),
    .A2(_09105_),
    .B1_N(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__and3b_1 _25769_ (.A_N(_09059_),
    .B(_09061_),
    .C(_09062_),
    .X(_09109_));
 sky130_fd_sc_hd__o21ai_4 _25770_ (.A1(_09104_),
    .A2(_09109_),
    .B1(_09102_),
    .Y(_09110_));
 sky130_fd_sc_hd__nand3b_4 _25771_ (.A_N(_09102_),
    .B(_09064_),
    .C(_09063_),
    .Y(_09111_));
 sky130_fd_sc_hd__nand3_4 _25772_ (.A(_09110_),
    .B(_09111_),
    .C(_09107_),
    .Y(_09112_));
 sky130_fd_sc_hd__a22oi_4 _25773_ (.A1(_09005_),
    .A2(_09006_),
    .B1(_09108_),
    .B2(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__a21oi_4 _25774_ (.A1(_09110_),
    .A2(_09111_),
    .B1(_09107_),
    .Y(_09114_));
 sky130_fd_sc_hd__nand2_4 _25775_ (.A(_09006_),
    .B(_09005_),
    .Y(_09115_));
 sky130_fd_sc_hd__nor3b_4 _25776_ (.A(_09114_),
    .B(_09115_),
    .C_N(_09112_),
    .Y(_09116_));
 sky130_fd_sc_hd__o21ai_4 _25777_ (.A1(_08926_),
    .A2(_08927_),
    .B1(_08924_),
    .Y(_09117_));
 sky130_fd_sc_hd__o21bai_4 _25778_ (.A1(_09113_),
    .A2(_09116_),
    .B1_N(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__nand3b_4 _25779_ (.A_N(_09115_),
    .B(_09108_),
    .C(_09112_),
    .Y(_09119_));
 sky130_fd_sc_hd__and3_1 _25780_ (.A(_09110_),
    .B(_09111_),
    .C(_09107_),
    .X(_09120_));
 sky130_fd_sc_hd__o21ai_2 _25781_ (.A1(_09114_),
    .A2(_09120_),
    .B1(_09115_),
    .Y(_09121_));
 sky130_fd_sc_hd__nand3_4 _25782_ (.A(_09119_),
    .B(_09121_),
    .C(_09117_),
    .Y(_09122_));
 sky130_fd_sc_hd__nor2_2 _25783_ (.A(_08797_),
    .B(_08812_),
    .Y(_09123_));
 sky130_fd_sc_hd__a21oi_4 _25784_ (.A1(_08811_),
    .A2(_08799_),
    .B1(_09123_),
    .Y(_09124_));
 sky130_fd_sc_hd__and2_1 _25785_ (.A(_08820_),
    .B(_08819_),
    .X(_09125_));
 sky130_fd_sc_hd__xor2_4 _25786_ (.A(_09124_),
    .B(_09125_),
    .X(_09126_));
 sky130_fd_sc_hd__a21oi_2 _25787_ (.A1(_09118_),
    .A2(_09122_),
    .B1(_09126_),
    .Y(_09127_));
 sky130_fd_sc_hd__nand3_4 _25788_ (.A(_09118_),
    .B(_09126_),
    .C(_09122_),
    .Y(_09128_));
 sky130_vsdinv _25789_ (.A(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__nand2_4 _25790_ (.A(_08940_),
    .B(_08933_),
    .Y(_09130_));
 sky130_fd_sc_hd__o21bai_4 _25791_ (.A1(_09127_),
    .A2(_09129_),
    .B1_N(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__a21o_1 _25792_ (.A1(_09118_),
    .A2(_09122_),
    .B1(_09126_),
    .X(_09132_));
 sky130_fd_sc_hd__nand3_4 _25793_ (.A(_09132_),
    .B(_09128_),
    .C(_09130_),
    .Y(_09133_));
 sky130_fd_sc_hd__nand2_1 _25794_ (.A(_09131_),
    .B(_09133_),
    .Y(_09134_));
 sky130_fd_sc_hd__a21boi_4 _25795_ (.A1(_08936_),
    .A2(_08617_),
    .B1_N(_08935_),
    .Y(_09135_));
 sky130_vsdinv _25796_ (.A(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__nand2_4 _25797_ (.A(_09134_),
    .B(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__nand3_4 _25798_ (.A(_09131_),
    .B(_09135_),
    .C(_09133_),
    .Y(_09138_));
 sky130_fd_sc_hd__nand2_2 _25799_ (.A(_08948_),
    .B(_08945_),
    .Y(_09139_));
 sky130_fd_sc_hd__a21oi_4 _25800_ (.A1(_09137_),
    .A2(_09138_),
    .B1(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__a21boi_2 _25801_ (.A1(_08943_),
    .A2(_08946_),
    .B1_N(_08945_),
    .Y(_09141_));
 sky130_fd_sc_hd__a21oi_4 _25802_ (.A1(_09131_),
    .A2(_09133_),
    .B1(_09135_),
    .Y(_09142_));
 sky130_fd_sc_hd__nor3b_4 _25803_ (.A(_09141_),
    .B(_09142_),
    .C_N(_09138_),
    .Y(_09143_));
 sky130_fd_sc_hd__nor2_4 _25804_ (.A(_09140_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__a21oi_2 _25805_ (.A1(_08955_),
    .A2(_08948_),
    .B1(_08952_),
    .Y(_09145_));
 sky130_fd_sc_hd__nor3_4 _25806_ (.A(_08950_),
    .B(_08947_),
    .C(_08949_),
    .Y(_09146_));
 sky130_fd_sc_hd__o21bai_1 _25807_ (.A1(_09145_),
    .A2(_08960_),
    .B1_N(_09146_),
    .Y(_09147_));
 sky130_fd_sc_hd__xor2_1 _25808_ (.A(_09144_),
    .B(_09147_),
    .X(_02654_));
 sky130_fd_sc_hd__o21a_2 _25809_ (.A1(_09011_),
    .A2(_09014_),
    .B1(_09012_),
    .X(_09148_));
 sky130_fd_sc_hd__a2bb2oi_4 _25810_ (.A1_N(_14418_),
    .A2_N(_09021_),
    .B1(_09020_),
    .B2(_09022_),
    .Y(_09149_));
 sky130_fd_sc_hd__nand2_4 _25811_ (.A(_07107_),
    .B(_05597_),
    .Y(_09150_));
 sky130_fd_sc_hd__or4_4 _25812_ (.A(_13985_),
    .B(_13990_),
    .C(_14394_),
    .D(_14400_),
    .X(_09151_));
 sky130_fd_sc_hd__buf_6 _25813_ (.A(_07264_),
    .X(_09152_));
 sky130_fd_sc_hd__buf_4 _25814_ (.A(_07102_),
    .X(_09153_));
 sky130_fd_sc_hd__a22o_1 _25815_ (.A1(_09152_),
    .A2(_05405_),
    .B1(_09153_),
    .B2(_05322_),
    .X(_09154_));
 sky130_fd_sc_hd__nand2_2 _25816_ (.A(_09151_),
    .B(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__xnor2_4 _25817_ (.A(_09150_),
    .B(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__xnor2_4 _25818_ (.A(_09149_),
    .B(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__xor2_4 _25819_ (.A(_09148_),
    .B(_09157_),
    .X(_09158_));
 sky130_fd_sc_hd__or2b_1 _25820_ (.A(_09032_),
    .B_N(_09027_),
    .X(_09159_));
 sky130_fd_sc_hd__o21ai_4 _25821_ (.A1(_09024_),
    .A2(_09033_),
    .B1(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__and2_2 _25822_ (.A(_07873_),
    .B(_05309_),
    .X(_09161_));
 sky130_fd_sc_hd__buf_4 _25823_ (.A(_13977_),
    .X(_09162_));
 sky130_fd_sc_hd__nand3_4 _25824_ (.A(_08396_),
    .B(_09162_),
    .C(_05819_),
    .Y(_09163_));
 sky130_fd_sc_hd__buf_2 _25825_ (.A(_13976_),
    .X(_09164_));
 sky130_fd_sc_hd__a22o_2 _25826_ (.A1(_08636_),
    .A2(_05819_),
    .B1(_09164_),
    .B2(_05875_),
    .X(_09165_));
 sky130_fd_sc_hd__o21ai_4 _25827_ (.A1(_14412_),
    .A2(_09163_),
    .B1(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__xor2_4 _25828_ (.A(_09161_),
    .B(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__buf_6 _25829_ (.A(_13966_),
    .X(_09168_));
 sky130_fd_sc_hd__buf_6 _25830_ (.A(_09025_),
    .X(_09169_));
 sky130_fd_sc_hd__nand3b_2 _25831_ (.A_N(_09029_),
    .B(_09169_),
    .C(_05178_),
    .Y(_09170_));
 sky130_fd_sc_hd__o31ai_4 _25832_ (.A1(_09168_),
    .A2(_14429_),
    .A3(_09031_),
    .B1(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__clkbuf_4 _25833_ (.A(\pcpi_mul.rs2[30] ),
    .X(_09172_));
 sky130_fd_sc_hd__and2_2 _25834_ (.A(_09172_),
    .B(_05091_),
    .X(_09173_));
 sky130_fd_sc_hd__clkbuf_4 _25835_ (.A(\pcpi_mul.rs2[31] ),
    .X(_09174_));
 sky130_fd_sc_hd__nand2_2 _25836_ (.A(_09174_),
    .B(_05959_),
    .Y(_09175_));
 sky130_fd_sc_hd__clkbuf_2 _25837_ (.A(\pcpi_mul.rs2[32] ),
    .X(_09176_));
 sky130_fd_sc_hd__and2b_1 _25838_ (.A_N(_04956_),
    .B(_09176_),
    .X(_09177_));
 sky130_fd_sc_hd__xor2_4 _25839_ (.A(_09175_),
    .B(_09177_),
    .X(_09178_));
 sky130_fd_sc_hd__xor2_4 _25840_ (.A(_09173_),
    .B(_09178_),
    .X(_09179_));
 sky130_fd_sc_hd__xor2_4 _25841_ (.A(_09171_),
    .B(_09179_),
    .X(_09180_));
 sky130_fd_sc_hd__xor2_4 _25842_ (.A(_09167_),
    .B(_09180_),
    .X(_09181_));
 sky130_fd_sc_hd__xnor2_4 _25843_ (.A(_09160_),
    .B(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__xnor2_4 _25844_ (.A(_09158_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__and2b_1 _25845_ (.A_N(_09035_),
    .B(_09017_),
    .X(_09184_));
 sky130_fd_sc_hd__a21o_2 _25846_ (.A1(_09034_),
    .A2(_09019_),
    .B1(_09184_),
    .X(_09185_));
 sky130_fd_sc_hd__nor2_2 _25847_ (.A(_09183_),
    .B(_09185_),
    .Y(_09186_));
 sky130_fd_sc_hd__nand2_4 _25848_ (.A(_09185_),
    .B(_09183_),
    .Y(_09187_));
 sky130_vsdinv _25849_ (.A(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__nor2_1 _25850_ (.A(_09046_),
    .B(_09052_),
    .Y(_09189_));
 sky130_fd_sc_hd__o21ba_2 _25851_ (.A1(_09045_),
    .A2(_09053_),
    .B1_N(_09189_),
    .X(_09190_));
 sky130_fd_sc_hd__and2_2 _25852_ (.A(_08261_),
    .B(_06279_),
    .X(_09191_));
 sky130_fd_sc_hd__nand3_4 _25853_ (.A(_08660_),
    .B(_08426_),
    .C(_06020_),
    .Y(_09192_));
 sky130_fd_sc_hd__a22o_2 _25854_ (.A1(_08662_),
    .A2(_06019_),
    .B1(_06896_),
    .B2(_06030_),
    .X(_09193_));
 sky130_fd_sc_hd__o21ai_4 _25855_ (.A1(_14360_),
    .A2(_09192_),
    .B1(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__xor2_4 _25856_ (.A(_09191_),
    .B(_09194_),
    .X(_09195_));
 sky130_fd_sc_hd__o21a_2 _25857_ (.A1(_06409_),
    .A2(_09048_),
    .B1(_09051_),
    .X(_09196_));
 sky130_fd_sc_hd__clkbuf_4 _25858_ (.A(_08269_),
    .X(_09197_));
 sky130_fd_sc_hd__buf_2 _25859_ (.A(_06412_),
    .X(_09198_));
 sky130_fd_sc_hd__a22o_1 _25860_ (.A1(_09197_),
    .A2(_06160_),
    .B1(_08668_),
    .B2(_09198_),
    .X(_09199_));
 sky130_fd_sc_hd__nand3_4 _25861_ (.A(_08269_),
    .B(_06647_),
    .C(_05512_),
    .Y(_09200_));
 sky130_fd_sc_hd__or2b_1 _25862_ (.A(_09200_),
    .B_N(_05611_),
    .X(_09201_));
 sky130_fd_sc_hd__o2bb2ai_1 _25863_ (.A1_N(_09199_),
    .A2_N(_09201_),
    .B1(_07123_),
    .B2(_14373_),
    .Y(_09202_));
 sky130_fd_sc_hd__o2111ai_4 _25864_ (.A1(_14378_),
    .A2(_09200_),
    .B1(_08673_),
    .C1(_05770_),
    .D1(_09199_),
    .Y(_09203_));
 sky130_fd_sc_hd__nand2_4 _25865_ (.A(_09202_),
    .B(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__xnor2_4 _25866_ (.A(_09196_),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__xor2_4 _25867_ (.A(_09195_),
    .B(_09205_),
    .X(_09206_));
 sky130_fd_sc_hd__nor2_1 _25868_ (.A(_09010_),
    .B(_09015_),
    .Y(_09207_));
 sky130_fd_sc_hd__o21bai_4 _25869_ (.A1(_09009_),
    .A2(_09016_),
    .B1_N(_09207_),
    .Y(_09208_));
 sky130_fd_sc_hd__xnor2_4 _25870_ (.A(_09206_),
    .B(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__xor2_4 _25871_ (.A(_09190_),
    .B(_09209_),
    .X(_09210_));
 sky130_fd_sc_hd__o21bai_4 _25872_ (.A1(_09186_),
    .A2(_09188_),
    .B1_N(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__nand3b_4 _25873_ (.A_N(_09186_),
    .B(_09210_),
    .C(_09187_),
    .Y(_09212_));
 sky130_fd_sc_hd__nand2_2 _25874_ (.A(_09061_),
    .B(_09037_),
    .Y(_09213_));
 sky130_fd_sc_hd__a21oi_4 _25875_ (.A1(_09211_),
    .A2(_09212_),
    .B1(_09213_),
    .Y(_09214_));
 sky130_vsdinv _25876_ (.A(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__nand3_4 _25877_ (.A(_09213_),
    .B(_09212_),
    .C(_09211_),
    .Y(_09216_));
 sky130_fd_sc_hd__or2b_1 _25878_ (.A(_09091_),
    .B_N(_09079_),
    .X(_09217_));
 sky130_fd_sc_hd__a21boi_4 _25879_ (.A1(_09090_),
    .A2(_09081_),
    .B1_N(_09217_),
    .Y(_09218_));
 sky130_fd_sc_hd__and2_1 _25880_ (.A(_09056_),
    .B(_09054_),
    .X(_09219_));
 sky130_fd_sc_hd__o21ba_2 _25881_ (.A1(_09040_),
    .A2(_09057_),
    .B1_N(_09219_),
    .X(_09220_));
 sky130_fd_sc_hd__and2_2 _25882_ (.A(_05206_),
    .B(_07769_),
    .X(_09221_));
 sky130_fd_sc_hd__clkbuf_8 _25883_ (.A(_14304_),
    .X(_09222_));
 sky130_fd_sc_hd__nand3_4 _25884_ (.A(_08333_),
    .B(_05274_),
    .C(_07575_),
    .Y(_09223_));
 sky130_fd_sc_hd__a22o_2 _25885_ (.A1(_08333_),
    .A2(_07575_),
    .B1(_05274_),
    .B2(_07775_),
    .X(_09224_));
 sky130_fd_sc_hd__o21ai_4 _25886_ (.A1(_09222_),
    .A2(_09223_),
    .B1(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__xnor2_4 _25887_ (.A(_09221_),
    .B(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__o21a_2 _25888_ (.A1(_14328_),
    .A2(_09073_),
    .B1(_09076_),
    .X(_09227_));
 sky130_fd_sc_hd__a22o_1 _25889_ (.A1(_14036_),
    .A2(\pcpi_mul.rs1[22] ),
    .B1(_05637_),
    .B2(_07204_),
    .X(_09228_));
 sky130_fd_sc_hd__nand3_4 _25890_ (.A(_05635_),
    .B(_05637_),
    .C(_14325_),
    .Y(_09229_));
 sky130_fd_sc_hd__or2b_1 _25891_ (.A(_09229_),
    .B_N(_07027_),
    .X(_09230_));
 sky130_fd_sc_hd__o2bb2ai_1 _25892_ (.A1_N(_09228_),
    .A2_N(_09230_),
    .B1(_14048_),
    .B2(_14315_),
    .Y(_09231_));
 sky130_fd_sc_hd__o2111ai_4 _25893_ (.A1(_14320_),
    .A2(_09229_),
    .B1(_05532_),
    .C1(_07038_),
    .D1(_09228_),
    .Y(_09232_));
 sky130_fd_sc_hd__nand2_4 _25894_ (.A(_09231_),
    .B(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__xnor2_4 _25895_ (.A(_09227_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__xnor2_4 _25896_ (.A(_09226_),
    .B(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__o21a_4 _25897_ (.A1(_09084_),
    .A2(_09087_),
    .B1(_09085_),
    .X(_09236_));
 sky130_fd_sc_hd__a2bb2oi_4 _25898_ (.A1_N(_14367_),
    .A2_N(_09042_),
    .B1(_09041_),
    .B2(_09043_),
    .Y(_09237_));
 sky130_fd_sc_hd__and2_2 _25899_ (.A(_05939_),
    .B(_06450_),
    .X(_09238_));
 sky130_fd_sc_hd__nand3_4 _25900_ (.A(_07294_),
    .B(_05814_),
    .C(_06431_),
    .Y(_09239_));
 sky130_fd_sc_hd__a22o_2 _25901_ (.A1(_05943_),
    .A2(_06583_),
    .B1(_05944_),
    .B2(_07746_),
    .X(_09240_));
 sky130_fd_sc_hd__o21ai_4 _25902_ (.A1(_14339_),
    .A2(_09239_),
    .B1(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__xor2_4 _25903_ (.A(_09238_),
    .B(_09241_),
    .X(_09242_));
 sky130_fd_sc_hd__xnor2_4 _25904_ (.A(_09237_),
    .B(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__xor2_4 _25905_ (.A(_09236_),
    .B(_09243_),
    .X(_09244_));
 sky130_fd_sc_hd__nor2_1 _25906_ (.A(_09083_),
    .B(_09088_),
    .Y(_09245_));
 sky130_fd_sc_hd__o21bai_4 _25907_ (.A1(_09082_),
    .A2(_09089_),
    .B1_N(_09245_),
    .Y(_09246_));
 sky130_fd_sc_hd__xnor2_4 _25908_ (.A(_09244_),
    .B(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__xnor2_4 _25909_ (.A(_09235_),
    .B(_09247_),
    .Y(_09248_));
 sky130_fd_sc_hd__xor2_4 _25910_ (.A(_09220_),
    .B(_09248_),
    .X(_09249_));
 sky130_fd_sc_hd__xnor2_2 _25911_ (.A(_09218_),
    .B(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__a21boi_1 _25912_ (.A1(_09215_),
    .A2(_09216_),
    .B1_N(_09250_),
    .Y(_09251_));
 sky130_fd_sc_hd__nand3b_4 _25913_ (.A_N(_09250_),
    .B(_09215_),
    .C(_09216_),
    .Y(_09252_));
 sky130_vsdinv _25914_ (.A(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__o21ai_4 _25915_ (.A1(_09102_),
    .A2(_09104_),
    .B1(_09064_),
    .Y(_09254_));
 sky130_fd_sc_hd__o21bai_2 _25916_ (.A1(_09251_),
    .A2(_09253_),
    .B1_N(_09254_),
    .Y(_09255_));
 sky130_fd_sc_hd__a21bo_2 _25917_ (.A1(_09215_),
    .A2(_09216_),
    .B1_N(_09250_),
    .X(_09256_));
 sky130_fd_sc_hd__nand3_4 _25918_ (.A(_09256_),
    .B(_09252_),
    .C(_09254_),
    .Y(_09257_));
 sky130_fd_sc_hd__nor2_1 _25919_ (.A(_08966_),
    .B(_08971_),
    .Y(_09258_));
 sky130_fd_sc_hd__o21ba_2 _25920_ (.A1(_08965_),
    .A2(_08972_),
    .B1_N(_09258_),
    .X(_09259_));
 sky130_fd_sc_hd__or2b_1 _25921_ (.A(_09078_),
    .B_N(_09069_),
    .X(_09260_));
 sky130_fd_sc_hd__o21ai_4 _25922_ (.A1(_09077_),
    .A2(_09070_),
    .B1(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__o21a_2 _25923_ (.A1(_08967_),
    .A2(_08970_),
    .B1(_08968_),
    .X(_09262_));
 sky130_fd_sc_hd__a2bb2oi_4 _25924_ (.A1_N(_14309_),
    .A2_N(_09066_),
    .B1(_09065_),
    .B2(_09067_),
    .Y(_09263_));
 sky130_fd_sc_hd__nand2_4 _25925_ (.A(_04998_),
    .B(_08806_),
    .Y(_09264_));
 sky130_fd_sc_hd__or4_4 _25926_ (.A(_14063_),
    .B(_14067_),
    .C(_14284_),
    .D(_14290_),
    .X(_09265_));
 sky130_fd_sc_hd__a22o_1 _25927_ (.A1(_05126_),
    .A2(_07584_),
    .B1(_05164_),
    .B2(_07784_),
    .X(_09266_));
 sky130_fd_sc_hd__nand2_2 _25928_ (.A(_09265_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__xnor2_4 _25929_ (.A(_09264_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__xnor2_4 _25930_ (.A(_09263_),
    .B(_09268_),
    .Y(_09269_));
 sky130_fd_sc_hd__xor2_4 _25931_ (.A(_09262_),
    .B(_09269_),
    .X(_09270_));
 sky130_fd_sc_hd__xnor2_4 _25932_ (.A(_09261_),
    .B(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__xor2_4 _25933_ (.A(_09259_),
    .B(_09271_),
    .X(_09272_));
 sky130_fd_sc_hd__and2_1 _25934_ (.A(_08973_),
    .B(_08964_),
    .X(_09273_));
 sky130_fd_sc_hd__o21ba_1 _25935_ (.A1(_08962_),
    .A2(_08974_),
    .B1_N(_09273_),
    .X(_09274_));
 sky130_fd_sc_hd__or2b_2 _25936_ (.A(_09272_),
    .B_N(_09274_),
    .X(_09275_));
 sky130_vsdinv _25937_ (.A(_09274_),
    .Y(_09276_));
 sky130_fd_sc_hd__nand2_2 _25938_ (.A(_09276_),
    .B(_09272_),
    .Y(_09277_));
 sky130_fd_sc_hd__o21a_4 _25939_ (.A1(_08985_),
    .A2(_08802_),
    .B1(_08981_),
    .X(_09278_));
 sky130_fd_sc_hd__buf_6 _25940_ (.A(_09278_),
    .X(_09279_));
 sky130_vsdinv _25941_ (.A(_08498_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand2_2 _25942_ (.A(_05117_),
    .B(_08171_),
    .Y(_09281_));
 sky130_fd_sc_hd__nand3b_4 _25943_ (.A_N(_09281_),
    .B(_12779_),
    .C(_08604_),
    .Y(_09282_));
 sky130_fd_sc_hd__clkbuf_4 _25944_ (.A(_12777_),
    .X(_09283_));
 sky130_fd_sc_hd__nand2_2 _25945_ (.A(_09283_),
    .B(_05515_),
    .Y(_09284_));
 sky130_fd_sc_hd__nand2_2 _25946_ (.A(_09281_),
    .B(_09284_),
    .Y(_09285_));
 sky130_fd_sc_hd__nand2_2 _25947_ (.A(_09282_),
    .B(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__xor2_4 _25948_ (.A(_09280_),
    .B(_09286_),
    .X(_09287_));
 sky130_fd_sc_hd__o21ai_4 _25949_ (.A1(_09280_),
    .A2(_08991_),
    .B1(_08989_),
    .Y(_09288_));
 sky130_fd_sc_hd__xnor2_4 _25950_ (.A(_09287_),
    .B(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__xor2_4 _25951_ (.A(_08986_),
    .B(_09289_),
    .X(_09290_));
 sky130_fd_sc_hd__or2_1 _25952_ (.A(_08988_),
    .B(_08992_),
    .X(_09291_));
 sky130_fd_sc_hd__o21a_2 _25953_ (.A1(_08987_),
    .A2(_08993_),
    .B1(_09291_),
    .X(_09292_));
 sky130_fd_sc_hd__xnor2_4 _25954_ (.A(_09290_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__xor2_4 _25955_ (.A(_09279_),
    .B(_09293_),
    .X(_09294_));
 sky130_fd_sc_hd__a21o_1 _25956_ (.A1(_09275_),
    .A2(_09277_),
    .B1(_09294_),
    .X(_09295_));
 sky130_fd_sc_hd__nand3_4 _25957_ (.A(_09275_),
    .B(_09294_),
    .C(_09277_),
    .Y(_09296_));
 sky130_fd_sc_hd__nand2_2 _25958_ (.A(_09101_),
    .B(_09096_),
    .Y(_09297_));
 sky130_fd_sc_hd__a21o_1 _25959_ (.A1(_09295_),
    .A2(_09296_),
    .B1(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__nand3_4 _25960_ (.A(_09297_),
    .B(_09295_),
    .C(_09296_),
    .Y(_09299_));
 sky130_fd_sc_hd__nand2_1 _25961_ (.A(_09298_),
    .B(_09299_),
    .Y(_09300_));
 sky130_fd_sc_hd__a21boi_1 _25962_ (.A1(_08978_),
    .A2(_08996_),
    .B1_N(_08980_),
    .Y(_09301_));
 sky130_fd_sc_hd__nand2_1 _25963_ (.A(_09300_),
    .B(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__nand3b_4 _25964_ (.A_N(_09301_),
    .B(_09298_),
    .C(_09299_),
    .Y(_09303_));
 sky130_fd_sc_hd__nand2_4 _25965_ (.A(_09302_),
    .B(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__a21boi_2 _25966_ (.A1(_09255_),
    .A2(_09257_),
    .B1_N(_09304_),
    .Y(_09305_));
 sky130_fd_sc_hd__a21oi_4 _25967_ (.A1(_09256_),
    .A2(_09252_),
    .B1(_09254_),
    .Y(_09306_));
 sky130_vsdinv _25968_ (.A(_09257_),
    .Y(_09307_));
 sky130_fd_sc_hd__nor3_4 _25969_ (.A(_09304_),
    .B(_09306_),
    .C(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__o21ai_2 _25970_ (.A1(_09114_),
    .A2(_09115_),
    .B1(_09112_),
    .Y(_09309_));
 sky130_fd_sc_hd__o21bai_4 _25971_ (.A1(_09305_),
    .A2(_09308_),
    .B1_N(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__o21ai_2 _25972_ (.A1(_09306_),
    .A2(_09307_),
    .B1(_09304_),
    .Y(_09311_));
 sky130_fd_sc_hd__nand3b_2 _25973_ (.A_N(_09304_),
    .B(_09255_),
    .C(_09257_),
    .Y(_09312_));
 sky130_fd_sc_hd__nand3_4 _25974_ (.A(_09311_),
    .B(_09309_),
    .C(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__nor2_2 _25975_ (.A(_08982_),
    .B(_08995_),
    .Y(_09314_));
 sky130_fd_sc_hd__a21oi_4 _25976_ (.A1(_08994_),
    .A2(_08984_),
    .B1(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__a21oi_4 _25977_ (.A1(_09005_),
    .A2(_09004_),
    .B1(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__and3_1 _25978_ (.A(_09005_),
    .B(_09004_),
    .C(_09315_),
    .X(_09317_));
 sky130_fd_sc_hd__nor2_4 _25979_ (.A(_09316_),
    .B(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__a21oi_2 _25980_ (.A1(_09310_),
    .A2(_09313_),
    .B1(_09318_),
    .Y(_09319_));
 sky130_fd_sc_hd__nand3_4 _25981_ (.A(_09310_),
    .B(_09318_),
    .C(_09313_),
    .Y(_09320_));
 sky130_vsdinv _25982_ (.A(_09320_),
    .Y(_09321_));
 sky130_vsdinv _25983_ (.A(_09126_),
    .Y(_09322_));
 sky130_fd_sc_hd__a21oi_2 _25984_ (.A1(_09119_),
    .A2(_09121_),
    .B1(_09117_),
    .Y(_09323_));
 sky130_fd_sc_hd__o21ai_4 _25985_ (.A1(_09322_),
    .A2(_09323_),
    .B1(_09122_),
    .Y(_09324_));
 sky130_fd_sc_hd__o21bai_4 _25986_ (.A1(_09319_),
    .A2(_09321_),
    .B1_N(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__o2bb2ai_2 _25987_ (.A1_N(_09313_),
    .A2_N(_09310_),
    .B1(_09316_),
    .B2(_09317_),
    .Y(_09326_));
 sky130_fd_sc_hd__nand3_4 _25988_ (.A(_09326_),
    .B(_09324_),
    .C(_09320_),
    .Y(_09327_));
 sky130_fd_sc_hd__a21oi_4 _25989_ (.A1(_08820_),
    .A2(_08819_),
    .B1(_09124_),
    .Y(_09328_));
 sky130_fd_sc_hd__a21oi_4 _25990_ (.A1(_09325_),
    .A2(_09327_),
    .B1(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__nand3_4 _25991_ (.A(_09325_),
    .B(_09328_),
    .C(_09327_),
    .Y(_09330_));
 sky130_vsdinv _25992_ (.A(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__a21oi_2 _25993_ (.A1(_09132_),
    .A2(_09128_),
    .B1(_09130_),
    .Y(_09332_));
 sky130_fd_sc_hd__o21ai_4 _25994_ (.A1(_09136_),
    .A2(_09332_),
    .B1(_09133_),
    .Y(_09333_));
 sky130_fd_sc_hd__o21bai_4 _25995_ (.A1(_09329_),
    .A2(_09331_),
    .B1_N(_09333_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand3b_4 _25996_ (.A_N(_09329_),
    .B(_09330_),
    .C(_09333_),
    .Y(_09335_));
 sky130_fd_sc_hd__nand2_8 _25997_ (.A(_09334_),
    .B(_09335_),
    .Y(_09336_));
 sky130_fd_sc_hd__nor3_4 _25998_ (.A(_09143_),
    .B(_09140_),
    .C(_08957_),
    .Y(_09337_));
 sky130_fd_sc_hd__nand3_2 _25999_ (.A(_09139_),
    .B(_09137_),
    .C(_09138_),
    .Y(_09338_));
 sky130_fd_sc_hd__o21ai_4 _26000_ (.A1(_08956_),
    .A2(_09140_),
    .B1(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__nand2_8 _26001_ (.A(_09337_),
    .B(_08958_),
    .Y(_09340_));
 sky130_fd_sc_hd__a31oi_4 _26002_ (.A1(_08554_),
    .A2(_08555_),
    .A3(_08566_),
    .B1(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__a211oi_4 _26003_ (.A1(_08959_),
    .A2(_09337_),
    .B1(_09339_),
    .C1(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__xor2_4 _26004_ (.A(_09336_),
    .B(net409),
    .X(_02655_));
 sky130_fd_sc_hd__nand2_2 _26005_ (.A(_09181_),
    .B(_09160_),
    .Y(_09343_));
 sky130_fd_sc_hd__or2b_2 _26006_ (.A(_09182_),
    .B_N(_09158_),
    .X(_09344_));
 sky130_fd_sc_hd__o21a_2 _26007_ (.A1(_09150_),
    .A2(_09155_),
    .B1(_09151_),
    .X(_09345_));
 sky130_fd_sc_hd__a2bb2oi_4 _26008_ (.A1_N(_14412_),
    .A2_N(_09163_),
    .B1(_09161_),
    .B2(_09165_),
    .Y(_09346_));
 sky130_fd_sc_hd__nand2_2 _26009_ (.A(_06888_),
    .B(_05604_),
    .Y(_09347_));
 sky130_fd_sc_hd__or4_4 _26010_ (.A(_13985_),
    .B(_13990_),
    .C(_14389_),
    .D(_14393_),
    .X(_09348_));
 sky130_fd_sc_hd__a22o_1 _26011_ (.A1(_08627_),
    .A2(_05322_),
    .B1(_08628_),
    .B2(_05424_),
    .X(_09349_));
 sky130_fd_sc_hd__nand2_2 _26012_ (.A(_09348_),
    .B(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__xnor2_4 _26013_ (.A(_09347_),
    .B(_09350_),
    .Y(_09351_));
 sky130_fd_sc_hd__xnor2_4 _26014_ (.A(_09346_),
    .B(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__xor2_4 _26015_ (.A(_09345_),
    .B(_09352_),
    .X(_09353_));
 sky130_fd_sc_hd__or2b_1 _26016_ (.A(_09179_),
    .B_N(_09171_),
    .X(_09354_));
 sky130_fd_sc_hd__o21ai_2 _26017_ (.A1(_09167_),
    .A2(_09180_),
    .B1(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__and2_2 _26018_ (.A(_08634_),
    .B(_05311_),
    .X(_09356_));
 sky130_fd_sc_hd__buf_4 _26019_ (.A(_13971_),
    .X(_09357_));
 sky130_fd_sc_hd__nand3_4 _26020_ (.A(_09357_),
    .B(_08637_),
    .C(_05875_),
    .Y(_09358_));
 sky130_fd_sc_hd__a22o_2 _26021_ (.A1(_08374_),
    .A2(_05228_),
    .B1(_09164_),
    .B2(_05309_),
    .X(_09359_));
 sky130_fd_sc_hd__o21ai_4 _26022_ (.A1(_14405_),
    .A2(_09358_),
    .B1(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__xor2_4 _26023_ (.A(_09356_),
    .B(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__nand3b_2 _26024_ (.A_N(_09175_),
    .B(_09169_),
    .C(_05580_),
    .Y(_09362_));
 sky130_fd_sc_hd__o31ai_4 _26025_ (.A1(_09168_),
    .A2(_14423_),
    .A3(_09178_),
    .B1(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__and2_2 _26026_ (.A(_08644_),
    .B(_05101_),
    .X(_09364_));
 sky130_fd_sc_hd__nand2_2 _26027_ (.A(_09174_),
    .B(_04983_),
    .Y(_09365_));
 sky130_fd_sc_hd__and2b_1 _26028_ (.A_N(_04960_),
    .B(_09176_),
    .X(_09366_));
 sky130_fd_sc_hd__xor2_4 _26029_ (.A(_09365_),
    .B(_09366_),
    .X(_09367_));
 sky130_fd_sc_hd__xor2_4 _26030_ (.A(_09364_),
    .B(_09367_),
    .X(_09368_));
 sky130_fd_sc_hd__xor2_4 _26031_ (.A(_09363_),
    .B(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__xor2_4 _26032_ (.A(_09361_),
    .B(_09369_),
    .X(_09370_));
 sky130_fd_sc_hd__xnor2_1 _26033_ (.A(_09355_),
    .B(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__xnor2_1 _26034_ (.A(_09353_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__a21bo_2 _26035_ (.A1(_09343_),
    .A2(_09344_),
    .B1_N(_09372_),
    .X(_09373_));
 sky130_fd_sc_hd__nand3b_4 _26036_ (.A_N(_09372_),
    .B(_09343_),
    .C(_09344_),
    .Y(_09374_));
 sky130_fd_sc_hd__nor2_1 _26037_ (.A(_09196_),
    .B(_09204_),
    .Y(_09375_));
 sky130_fd_sc_hd__o21ba_2 _26038_ (.A1(_09195_),
    .A2(_09205_),
    .B1_N(_09375_),
    .X(_09376_));
 sky130_fd_sc_hd__and2_2 _26039_ (.A(_06346_),
    .B(_08342_),
    .X(_09377_));
 sky130_fd_sc_hd__nand3_4 _26040_ (.A(_08422_),
    .B(_08859_),
    .C(_06147_),
    .Y(_09378_));
 sky130_fd_sc_hd__buf_6 _26041_ (.A(_06185_),
    .X(_09379_));
 sky130_fd_sc_hd__a22o_2 _26042_ (.A1(_08662_),
    .A2(_06285_),
    .B1(_09379_),
    .B2(_06438_),
    .X(_09380_));
 sky130_fd_sc_hd__o21ai_4 _26043_ (.A1(_14354_),
    .A2(_09378_),
    .B1(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__xor2_4 _26044_ (.A(_09377_),
    .B(_09381_),
    .X(_09382_));
 sky130_fd_sc_hd__o21a_2 _26045_ (.A1(_14379_),
    .A2(_09200_),
    .B1(_09203_),
    .X(_09383_));
 sky130_fd_sc_hd__a22o_1 _26046_ (.A1(_09197_),
    .A2(_05691_),
    .B1(_08668_),
    .B2(_05905_),
    .X(_09384_));
 sky130_fd_sc_hd__nand3_4 _26047_ (.A(_08431_),
    .B(_08432_),
    .C(_09198_),
    .Y(_09385_));
 sky130_fd_sc_hd__or2b_1 _26048_ (.A(_09385_),
    .B_N(_05700_),
    .X(_09386_));
 sky130_fd_sc_hd__o2bb2ai_1 _26049_ (.A1_N(_09384_),
    .A2_N(_09386_),
    .B1(_14006_),
    .B2(_14367_),
    .Y(_09387_));
 sky130_fd_sc_hd__buf_6 _26050_ (.A(_06649_),
    .X(_09388_));
 sky130_fd_sc_hd__o2111ai_4 _26051_ (.A1(_14372_),
    .A2(_09385_),
    .B1(_09388_),
    .C1(_06020_),
    .D1(_09384_),
    .Y(_09389_));
 sky130_fd_sc_hd__nand2_4 _26052_ (.A(_09387_),
    .B(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__xnor2_4 _26053_ (.A(_09383_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__xor2_4 _26054_ (.A(_09382_),
    .B(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__nor2_1 _26055_ (.A(_09149_),
    .B(_09156_),
    .Y(_09393_));
 sky130_fd_sc_hd__o21bai_4 _26056_ (.A1(_09148_),
    .A2(_09157_),
    .B1_N(_09393_),
    .Y(_09394_));
 sky130_fd_sc_hd__xnor2_4 _26057_ (.A(_09392_),
    .B(_09394_),
    .Y(_09395_));
 sky130_fd_sc_hd__xor2_4 _26058_ (.A(_09376_),
    .B(_09395_),
    .X(_09396_));
 sky130_fd_sc_hd__a21oi_2 _26059_ (.A1(_09373_),
    .A2(_09374_),
    .B1(_09396_),
    .Y(_09397_));
 sky130_vsdinv _26060_ (.A(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__nand3_4 _26061_ (.A(_09373_),
    .B(_09396_),
    .C(_09374_),
    .Y(_09399_));
 sky130_fd_sc_hd__nand2_4 _26062_ (.A(_09212_),
    .B(_09187_),
    .Y(_09400_));
 sky130_fd_sc_hd__a21o_1 _26063_ (.A1(_09398_),
    .A2(_09399_),
    .B1(_09400_),
    .X(_09401_));
 sky130_fd_sc_hd__nand3b_4 _26064_ (.A_N(_09397_),
    .B(_09400_),
    .C(_09399_),
    .Y(_09402_));
 sky130_fd_sc_hd__nand2_1 _26065_ (.A(_09246_),
    .B(_09244_),
    .Y(_09403_));
 sky130_fd_sc_hd__or2b_1 _26066_ (.A(_09247_),
    .B_N(_09235_),
    .X(_09404_));
 sky130_fd_sc_hd__and2_2 _26067_ (.A(_05205_),
    .B(_08779_),
    .X(_09405_));
 sky130_fd_sc_hd__nand3_4 _26068_ (.A(_05359_),
    .B(_05363_),
    .C(_07568_),
    .Y(_09406_));
 sky130_fd_sc_hd__a22o_1 _26069_ (.A1(_05361_),
    .A2(_07216_),
    .B1(_05363_),
    .B2(_08782_),
    .X(_09407_));
 sky130_fd_sc_hd__o21ai_2 _26070_ (.A1(_14297_),
    .A2(_09406_),
    .B1(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__xnor2_2 _26071_ (.A(_09405_),
    .B(_09408_),
    .Y(_09409_));
 sky130_fd_sc_hd__o21a_2 _26072_ (.A1(_14320_),
    .A2(_09229_),
    .B1(_09232_),
    .X(_09410_));
 sky130_fd_sc_hd__a22o_1 _26073_ (.A1(_05635_),
    .A2(_07204_),
    .B1(_05637_),
    .B2(_06956_),
    .X(_09411_));
 sky130_fd_sc_hd__nand3_4 _26074_ (.A(_05730_),
    .B(_05732_),
    .C(\pcpi_mul.rs1[23] ),
    .Y(_09412_));
 sky130_fd_sc_hd__or2b_1 _26075_ (.A(_09412_),
    .B_N(_07038_),
    .X(_09413_));
 sky130_fd_sc_hd__o2bb2ai_1 _26076_ (.A1_N(_09411_),
    .A2_N(_09413_),
    .B1(_14046_),
    .B2(_14308_),
    .Y(_09414_));
 sky130_fd_sc_hd__o2111ai_4 _26077_ (.A1(_14313_),
    .A2(_09412_),
    .B1(_05532_),
    .C1(_07209_),
    .D1(_09411_),
    .Y(_09415_));
 sky130_fd_sc_hd__nand2_4 _26078_ (.A(_09414_),
    .B(_09415_),
    .Y(_09416_));
 sky130_fd_sc_hd__xnor2_2 _26079_ (.A(_09410_),
    .B(_09416_),
    .Y(_09417_));
 sky130_fd_sc_hd__xnor2_2 _26080_ (.A(_09409_),
    .B(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__nor2_1 _26081_ (.A(_09237_),
    .B(_09242_),
    .Y(_09419_));
 sky130_fd_sc_hd__o21bai_4 _26082_ (.A1(_09236_),
    .A2(_09243_),
    .B1_N(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__a2bb2oi_4 _26083_ (.A1_N(_14342_),
    .A2_N(_09239_),
    .B1(_09238_),
    .B2(_09240_),
    .Y(_09421_));
 sky130_fd_sc_hd__a2bb2oi_4 _26084_ (.A1_N(_14360_),
    .A2_N(_09192_),
    .B1(_09191_),
    .B2(_09193_),
    .Y(_09422_));
 sky130_fd_sc_hd__and2_2 _26085_ (.A(_05717_),
    .B(_07033_),
    .X(_09423_));
 sky130_fd_sc_hd__nand3_4 _26086_ (.A(_05943_),
    .B(_06071_),
    .C(_07046_),
    .Y(_09424_));
 sky130_fd_sc_hd__a22o_2 _26087_ (.A1(_08354_),
    .A2(_06296_),
    .B1(_08355_),
    .B2(_07048_),
    .X(_09425_));
 sky130_fd_sc_hd__o21ai_4 _26088_ (.A1(_14333_),
    .A2(_09424_),
    .B1(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__xor2_4 _26089_ (.A(_09423_),
    .B(_09426_),
    .X(_09427_));
 sky130_fd_sc_hd__xnor2_4 _26090_ (.A(_09422_),
    .B(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__xor2_4 _26091_ (.A(_09421_),
    .B(_09428_),
    .X(_09429_));
 sky130_fd_sc_hd__xnor2_1 _26092_ (.A(_09420_),
    .B(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__xnor2_1 _26093_ (.A(_09418_),
    .B(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__and2_1 _26094_ (.A(_09208_),
    .B(_09206_),
    .X(_09432_));
 sky130_fd_sc_hd__o21ba_1 _26095_ (.A1(_09190_),
    .A2(_09209_),
    .B1_N(_09432_),
    .X(_09433_));
 sky130_fd_sc_hd__xor2_1 _26096_ (.A(_09431_),
    .B(_09433_),
    .X(_09434_));
 sky130_fd_sc_hd__a21o_1 _26097_ (.A1(_09403_),
    .A2(_09404_),
    .B1(_09434_),
    .X(_09435_));
 sky130_fd_sc_hd__nand3_1 _26098_ (.A(_09434_),
    .B(_09403_),
    .C(_09404_),
    .Y(_09436_));
 sky130_fd_sc_hd__nand2_2 _26099_ (.A(_09435_),
    .B(_09436_),
    .Y(_09437_));
 sky130_vsdinv _26100_ (.A(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__a21oi_1 _26101_ (.A1(_09401_),
    .A2(_09402_),
    .B1(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__nand3_4 _26102_ (.A(_09401_),
    .B(_09438_),
    .C(_09402_),
    .Y(_09440_));
 sky130_vsdinv _26103_ (.A(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__o21ai_4 _26104_ (.A1(_09214_),
    .A2(_09250_),
    .B1(_09216_),
    .Y(_09442_));
 sky130_fd_sc_hd__o21bai_2 _26105_ (.A1(_09439_),
    .A2(_09441_),
    .B1_N(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__a21o_1 _26106_ (.A1(_09401_),
    .A2(_09402_),
    .B1(_09438_),
    .X(_09444_));
 sky130_fd_sc_hd__nand3_4 _26107_ (.A(_09444_),
    .B(_09440_),
    .C(_09442_),
    .Y(_09445_));
 sky130_fd_sc_hd__nand2_1 _26108_ (.A(_09443_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__nor2_2 _26109_ (.A(_09259_),
    .B(_09271_),
    .Y(_09447_));
 sky130_fd_sc_hd__a21oi_4 _26110_ (.A1(_09261_),
    .A2(_09270_),
    .B1(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__nor2_1 _26111_ (.A(_09263_),
    .B(_09268_),
    .Y(_09449_));
 sky130_fd_sc_hd__o21ba_2 _26112_ (.A1(_09262_),
    .A2(_09269_),
    .B1_N(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__or2b_1 _26113_ (.A(_09234_),
    .B_N(_09226_),
    .X(_09451_));
 sky130_fd_sc_hd__o21ai_4 _26114_ (.A1(_09233_),
    .A2(_09227_),
    .B1(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__o21a_2 _26115_ (.A1(_09264_),
    .A2(_09267_),
    .B1(_09265_),
    .X(_09453_));
 sky130_fd_sc_hd__a2bb2oi_4 _26116_ (.A1_N(_09222_),
    .A2_N(_09223_),
    .B1(_09221_),
    .B2(_09224_),
    .Y(_09454_));
 sky130_fd_sc_hd__nand2_4 _26117_ (.A(_04999_),
    .B(_08492_),
    .Y(_09455_));
 sky130_fd_sc_hd__or4_4 _26118_ (.A(_14063_),
    .B(_14067_),
    .C(_14278_),
    .D(_14285_),
    .X(_09456_));
 sky130_fd_sc_hd__a22o_1 _26119_ (.A1(_05132_),
    .A2(_08487_),
    .B1(_05065_),
    .B2(_08165_),
    .X(_09457_));
 sky130_fd_sc_hd__nand2_2 _26120_ (.A(_09456_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__xnor2_4 _26121_ (.A(_09455_),
    .B(_09458_),
    .Y(_09459_));
 sky130_fd_sc_hd__xnor2_4 _26122_ (.A(_09454_),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__xor2_4 _26123_ (.A(_09453_),
    .B(_09460_),
    .X(_09461_));
 sky130_fd_sc_hd__xnor2_4 _26124_ (.A(_09452_),
    .B(_09461_),
    .Y(_09462_));
 sky130_fd_sc_hd__xor2_1 _26125_ (.A(_09450_),
    .B(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__or2b_2 _26126_ (.A(_09448_),
    .B_N(_09463_),
    .X(_09464_));
 sky130_fd_sc_hd__nor2_2 _26127_ (.A(_09450_),
    .B(_09462_),
    .Y(_09465_));
 sky130_fd_sc_hd__and2_1 _26128_ (.A(_09462_),
    .B(_09450_),
    .X(_09466_));
 sky130_fd_sc_hd__o21ai_2 _26129_ (.A1(_09465_),
    .A2(_09466_),
    .B1(_09448_),
    .Y(_09467_));
 sky130_fd_sc_hd__buf_6 _26130_ (.A(_12779_),
    .X(_09468_));
 sky130_fd_sc_hd__o21a_2 _26131_ (.A1(_05316_),
    .A2(_08604_),
    .B1(_09468_),
    .X(_09469_));
 sky130_fd_sc_hd__o21a_2 _26132_ (.A1(_14075_),
    .A2(_09284_),
    .B1(_09469_),
    .X(_09470_));
 sky130_fd_sc_hd__a22oi_4 _26133_ (.A1(_04714_),
    .A2(_09285_),
    .B1(_09282_),
    .B2(_09280_),
    .Y(_09471_));
 sky130_fd_sc_hd__xor2_4 _26134_ (.A(_09470_),
    .B(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__xor2_4 _26135_ (.A(_08986_),
    .B(_09472_),
    .X(_09473_));
 sky130_fd_sc_hd__and2_1 _26136_ (.A(_09288_),
    .B(_09287_),
    .X(_09474_));
 sky130_fd_sc_hd__o21bai_4 _26137_ (.A1(_08987_),
    .A2(_09289_),
    .B1_N(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__xnor2_4 _26138_ (.A(_09473_),
    .B(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__xor2_4 _26139_ (.A(_09279_),
    .B(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__a21o_1 _26140_ (.A1(_09464_),
    .A2(_09467_),
    .B1(_09477_),
    .X(_09478_));
 sky130_fd_sc_hd__nand3_4 _26141_ (.A(_09464_),
    .B(_09467_),
    .C(_09477_),
    .Y(_09479_));
 sky130_fd_sc_hd__and2b_1 _26142_ (.A_N(_09220_),
    .B(_09248_),
    .X(_09480_));
 sky130_fd_sc_hd__o21bai_4 _26143_ (.A1(_09218_),
    .A2(_09249_),
    .B1_N(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__a21o_2 _26144_ (.A1(_09478_),
    .A2(_09479_),
    .B1(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__nand3_4 _26145_ (.A(_09478_),
    .B(_09481_),
    .C(_09479_),
    .Y(_09483_));
 sky130_vsdinv _26146_ (.A(_09277_),
    .Y(_09484_));
 sky130_fd_sc_hd__a21oi_1 _26147_ (.A1(_09275_),
    .A2(_09294_),
    .B1(_09484_),
    .Y(_09485_));
 sky130_vsdinv _26148_ (.A(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__a21o_1 _26149_ (.A1(_09482_),
    .A2(_09483_),
    .B1(_09486_),
    .X(_09487_));
 sky130_fd_sc_hd__nand3_4 _26150_ (.A(_09482_),
    .B(_09486_),
    .C(_09483_),
    .Y(_09488_));
 sky130_fd_sc_hd__nand2_2 _26151_ (.A(_09487_),
    .B(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__nand2_2 _26152_ (.A(_09446_),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__nand3b_4 _26153_ (.A_N(_09489_),
    .B(_09443_),
    .C(_09445_),
    .Y(_09491_));
 sky130_fd_sc_hd__o21ai_4 _26154_ (.A1(_09304_),
    .A2(_09306_),
    .B1(_09257_),
    .Y(_09492_));
 sky130_fd_sc_hd__a21o_1 _26155_ (.A1(_09490_),
    .A2(_09491_),
    .B1(_09492_),
    .X(_09493_));
 sky130_fd_sc_hd__nand3_4 _26156_ (.A(_09490_),
    .B(_09491_),
    .C(_09492_),
    .Y(_09494_));
 sky130_fd_sc_hd__nor2_1 _26157_ (.A(_09290_),
    .B(_09292_),
    .Y(_09495_));
 sky130_fd_sc_hd__o21bai_4 _26158_ (.A1(_09279_),
    .A2(_09293_),
    .B1_N(_09495_),
    .Y(_09496_));
 sky130_fd_sc_hd__nand2_2 _26159_ (.A(_09303_),
    .B(_09299_),
    .Y(_09497_));
 sky130_fd_sc_hd__xor2_4 _26160_ (.A(_09496_),
    .B(_09497_),
    .X(_09498_));
 sky130_fd_sc_hd__a21oi_1 _26161_ (.A1(_09493_),
    .A2(_09494_),
    .B1(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__nand3_4 _26162_ (.A(_09493_),
    .B(_09498_),
    .C(_09494_),
    .Y(_09500_));
 sky130_vsdinv _26163_ (.A(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__nand2_4 _26164_ (.A(_09320_),
    .B(_09313_),
    .Y(_09502_));
 sky130_fd_sc_hd__o21bai_2 _26165_ (.A1(_09499_),
    .A2(_09501_),
    .B1_N(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__a21oi_4 _26166_ (.A1(_09490_),
    .A2(_09491_),
    .B1(_09492_),
    .Y(_09504_));
 sky130_vsdinv _26167_ (.A(_09494_),
    .Y(_09505_));
 sky130_fd_sc_hd__o21bai_4 _26168_ (.A1(_09504_),
    .A2(_09505_),
    .B1_N(_09498_),
    .Y(_09506_));
 sky130_fd_sc_hd__nand3_4 _26169_ (.A(_09502_),
    .B(_09506_),
    .C(_09500_),
    .Y(_09507_));
 sky130_fd_sc_hd__a21oi_1 _26170_ (.A1(_09503_),
    .A2(_09507_),
    .B1(_09316_),
    .Y(_09508_));
 sky130_vsdinv _26171_ (.A(_09316_),
    .Y(_09509_));
 sky130_fd_sc_hd__a21oi_4 _26172_ (.A1(_09506_),
    .A2(_09500_),
    .B1(_09502_),
    .Y(_09510_));
 sky130_fd_sc_hd__nor3b_4 _26173_ (.A(_09509_),
    .B(_09510_),
    .C_N(_09507_),
    .Y(_09511_));
 sky130_fd_sc_hd__nand2_2 _26174_ (.A(_09330_),
    .B(_09327_),
    .Y(_09512_));
 sky130_fd_sc_hd__o21bai_2 _26175_ (.A1(_09508_),
    .A2(_09511_),
    .B1_N(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__a21boi_1 _26176_ (.A1(_09001_),
    .A2(_09003_),
    .B1_N(_09004_),
    .Y(_09514_));
 sky130_fd_sc_hd__o2bb2ai_1 _26177_ (.A1_N(_09507_),
    .A2_N(_09503_),
    .B1(_09514_),
    .B2(_09315_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand3_2 _26178_ (.A(_09503_),
    .B(_09316_),
    .C(_09507_),
    .Y(_09516_));
 sky130_fd_sc_hd__nand3_4 _26179_ (.A(_09515_),
    .B(_09512_),
    .C(_09516_),
    .Y(_09517_));
 sky130_fd_sc_hd__nand2_4 _26180_ (.A(_09513_),
    .B(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__o21ai_4 _26181_ (.A1(_09336_),
    .A2(net409),
    .B1(_09335_),
    .Y(_09519_));
 sky130_fd_sc_hd__xnor2_4 _26182_ (.A(_09518_),
    .B(_09519_),
    .Y(_02656_));
 sky130_fd_sc_hd__o21a_2 _26183_ (.A1(_09347_),
    .A2(_09350_),
    .B1(_09348_),
    .X(_09520_));
 sky130_fd_sc_hd__a2bb2oi_4 _26184_ (.A1_N(_14406_),
    .A2_N(_09358_),
    .B1(_09356_),
    .B2(_09359_),
    .Y(_09521_));
 sky130_fd_sc_hd__nand2_2 _26185_ (.A(_06888_),
    .B(_05692_),
    .Y(_09522_));
 sky130_fd_sc_hd__or4_4 _26186_ (.A(_13985_),
    .B(_13990_),
    .C(_14383_),
    .D(_14388_),
    .X(_09523_));
 sky130_fd_sc_hd__a22o_1 _26187_ (.A1(_08404_),
    .A2(_08264_),
    .B1(_08628_),
    .B2(_06160_),
    .X(_09524_));
 sky130_fd_sc_hd__nand2_2 _26188_ (.A(_09523_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__xnor2_2 _26189_ (.A(_09522_),
    .B(_09525_),
    .Y(_09526_));
 sky130_fd_sc_hd__xnor2_2 _26190_ (.A(_09521_),
    .B(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__xor2_2 _26191_ (.A(_09520_),
    .B(_09527_),
    .X(_09528_));
 sky130_fd_sc_hd__or2b_1 _26192_ (.A(_09368_),
    .B_N(_09363_),
    .X(_09529_));
 sky130_fd_sc_hd__o21ai_2 _26193_ (.A1(_09361_),
    .A2(_09369_),
    .B1(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__and2_2 _26194_ (.A(_08634_),
    .B(_05414_),
    .X(_09531_));
 sky130_fd_sc_hd__nand3_4 _26195_ (.A(_09357_),
    .B(_09162_),
    .C(_05309_),
    .Y(_09532_));
 sky130_fd_sc_hd__a22o_2 _26196_ (.A1(_08636_),
    .A2(_05237_),
    .B1(_09164_),
    .B2(_05311_),
    .X(_09533_));
 sky130_fd_sc_hd__o21ai_4 _26197_ (.A1(_05874_),
    .A2(_09532_),
    .B1(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__xor2_4 _26198_ (.A(_09531_),
    .B(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__nand3b_2 _26199_ (.A_N(_09365_),
    .B(_09169_),
    .C(_05247_),
    .Y(_09536_));
 sky130_fd_sc_hd__o31ai_4 _26200_ (.A1(_09168_),
    .A2(_14418_),
    .A3(_09367_),
    .B1(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__and2_2 _26201_ (.A(_09172_),
    .B(_05106_),
    .X(_09538_));
 sky130_fd_sc_hd__nand2_2 _26202_ (.A(_08646_),
    .B(_05047_),
    .Y(_09539_));
 sky130_fd_sc_hd__and2b_1 _26203_ (.A_N(_05098_),
    .B(_08383_),
    .X(_09540_));
 sky130_fd_sc_hd__xor2_4 _26204_ (.A(_09539_),
    .B(_09540_),
    .X(_09541_));
 sky130_fd_sc_hd__xor2_4 _26205_ (.A(_09538_),
    .B(_09541_),
    .X(_09542_));
 sky130_fd_sc_hd__xor2_4 _26206_ (.A(_09537_),
    .B(_09542_),
    .X(_09543_));
 sky130_fd_sc_hd__xor2_4 _26207_ (.A(_09535_),
    .B(_09543_),
    .X(_09544_));
 sky130_fd_sc_hd__xnor2_1 _26208_ (.A(_09530_),
    .B(_09544_),
    .Y(_09545_));
 sky130_fd_sc_hd__xnor2_1 _26209_ (.A(_09528_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__or2_1 _26210_ (.A(_09355_),
    .B(_09370_),
    .X(_09547_));
 sky130_fd_sc_hd__nand2_1 _26211_ (.A(_09370_),
    .B(_09355_),
    .Y(_09548_));
 sky130_fd_sc_hd__a21boi_4 _26212_ (.A1(_09547_),
    .A2(_09353_),
    .B1_N(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__or2b_2 _26213_ (.A(_09546_),
    .B_N(_09549_),
    .X(_09550_));
 sky130_fd_sc_hd__or2b_2 _26214_ (.A(_09549_),
    .B_N(_09546_),
    .X(_09551_));
 sky130_fd_sc_hd__nor2_1 _26215_ (.A(_09383_),
    .B(_09390_),
    .Y(_09552_));
 sky130_fd_sc_hd__o21ba_4 _26216_ (.A1(_09382_),
    .A2(_09391_),
    .B1_N(_09552_),
    .X(_09553_));
 sky130_fd_sc_hd__nor2_1 _26217_ (.A(_09346_),
    .B(_09351_),
    .Y(_09554_));
 sky130_fd_sc_hd__o21bai_4 _26218_ (.A1(_09345_),
    .A2(_09352_),
    .B1_N(_09554_),
    .Y(_09555_));
 sky130_fd_sc_hd__and2_2 _26219_ (.A(_06346_),
    .B(_06441_),
    .X(_09556_));
 sky130_fd_sc_hd__nand3_4 _26220_ (.A(_08422_),
    .B(_08859_),
    .C(_06438_),
    .Y(_09557_));
 sky130_fd_sc_hd__a22o_2 _26221_ (.A1(_08425_),
    .A2(_06279_),
    .B1(_09379_),
    .B2(_08342_),
    .X(_09558_));
 sky130_fd_sc_hd__o21ai_4 _26222_ (.A1(_14347_),
    .A2(_09557_),
    .B1(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__xor2_4 _26223_ (.A(_09556_),
    .B(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__o21a_2 _26224_ (.A1(_14373_),
    .A2(_09385_),
    .B1(_09389_),
    .X(_09561_));
 sky130_fd_sc_hd__nand2_4 _26225_ (.A(_08673_),
    .B(_06147_),
    .Y(_09562_));
 sky130_fd_sc_hd__or4_4 _26226_ (.A(_13999_),
    .B(_14002_),
    .C(_14365_),
    .D(_14371_),
    .X(_09563_));
 sky130_fd_sc_hd__a22o_1 _26227_ (.A1(_09197_),
    .A2(_05769_),
    .B1(_08668_),
    .B2(_08720_),
    .X(_09564_));
 sky130_fd_sc_hd__nand2_2 _26228_ (.A(_09563_),
    .B(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__xnor2_4 _26229_ (.A(_09562_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__xnor2_4 _26230_ (.A(_09561_),
    .B(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__xor2_4 _26231_ (.A(_09560_),
    .B(_09567_),
    .X(_09568_));
 sky130_fd_sc_hd__xnor2_4 _26232_ (.A(_09555_),
    .B(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__xor2_4 _26233_ (.A(_09553_),
    .B(_09569_),
    .X(_09570_));
 sky130_fd_sc_hd__a21o_1 _26234_ (.A1(_09550_),
    .A2(_09551_),
    .B1(_09570_),
    .X(_09571_));
 sky130_fd_sc_hd__nand3_4 _26235_ (.A(_09570_),
    .B(_09550_),
    .C(_09551_),
    .Y(_09572_));
 sky130_fd_sc_hd__nand2_2 _26236_ (.A(_09399_),
    .B(_09373_),
    .Y(_09573_));
 sky130_fd_sc_hd__a21o_2 _26237_ (.A1(_09571_),
    .A2(_09572_),
    .B1(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__nand3_4 _26238_ (.A(_09573_),
    .B(_09572_),
    .C(_09571_),
    .Y(_09575_));
 sky130_fd_sc_hd__or2b_1 _26239_ (.A(_09430_),
    .B_N(_09418_),
    .X(_09576_));
 sky130_fd_sc_hd__a21boi_4 _26240_ (.A1(_09429_),
    .A2(_09420_),
    .B1_N(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__and2_2 _26241_ (.A(_05205_),
    .B(_07784_),
    .X(_09578_));
 sky130_fd_sc_hd__nand3_4 _26242_ (.A(_05582_),
    .B(_05273_),
    .C(_07485_),
    .Y(_09579_));
 sky130_fd_sc_hd__a22o_2 _26243_ (.A1(_05361_),
    .A2(_08782_),
    .B1(_05363_),
    .B2(_08779_),
    .X(_09580_));
 sky130_fd_sc_hd__o21ai_4 _26244_ (.A1(_14291_),
    .A2(_09579_),
    .B1(_09580_),
    .Y(_09581_));
 sky130_fd_sc_hd__xnor2_4 _26245_ (.A(_09578_),
    .B(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__o21a_4 _26246_ (.A1(_14314_),
    .A2(_09412_),
    .B1(_09415_),
    .X(_09583_));
 sky130_fd_sc_hd__a22o_1 _26247_ (.A1(_05635_),
    .A2(_06956_),
    .B1(_08199_),
    .B2(_07786_),
    .X(_09584_));
 sky130_fd_sc_hd__nand3_4 _26248_ (.A(_14036_),
    .B(_05732_),
    .C(\pcpi_mul.rs1[24] ),
    .Y(_09585_));
 sky130_fd_sc_hd__or2b_1 _26249_ (.A(_09585_),
    .B_N(_07786_),
    .X(_09586_));
 sky130_fd_sc_hd__o2bb2ai_1 _26250_ (.A1_N(_09584_),
    .A2_N(_09586_),
    .B1(_06207_),
    .B2(_14303_),
    .Y(_09587_));
 sky130_fd_sc_hd__o2111ai_4 _26251_ (.A1(_14307_),
    .A2(_09585_),
    .B1(_05441_),
    .C1(_07216_),
    .D1(_09584_),
    .Y(_09588_));
 sky130_fd_sc_hd__nand2_4 _26252_ (.A(_09587_),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__xnor2_4 _26253_ (.A(_09583_),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__xnor2_4 _26254_ (.A(_09582_),
    .B(_09590_),
    .Y(_09591_));
 sky130_fd_sc_hd__nor2_1 _26255_ (.A(_09422_),
    .B(_09427_),
    .Y(_09592_));
 sky130_fd_sc_hd__o21bai_4 _26256_ (.A1(_09421_),
    .A2(_09428_),
    .B1_N(_09592_),
    .Y(_09593_));
 sky130_fd_sc_hd__a2bb2oi_4 _26257_ (.A1_N(_14335_),
    .A2_N(_09424_),
    .B1(_09423_),
    .B2(_09425_),
    .Y(_09594_));
 sky130_fd_sc_hd__a2bb2oi_4 _26258_ (.A1_N(_08338_),
    .A2_N(_09378_),
    .B1(_09377_),
    .B2(_09380_),
    .Y(_09595_));
 sky130_fd_sc_hd__and2_2 _26259_ (.A(_05717_),
    .B(_07036_),
    .X(_09596_));
 sky130_fd_sc_hd__nand3_4 _26260_ (.A(_05941_),
    .B(_05814_),
    .C(_06760_),
    .Y(_09597_));
 sky130_fd_sc_hd__a22o_2 _26261_ (.A1(_06067_),
    .A2(_07048_),
    .B1(_06071_),
    .B2(_06939_),
    .X(_09598_));
 sky130_fd_sc_hd__o21ai_4 _26262_ (.A1(_14327_),
    .A2(_09597_),
    .B1(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__xor2_4 _26263_ (.A(_09596_),
    .B(_09599_),
    .X(_09600_));
 sky130_fd_sc_hd__xnor2_4 _26264_ (.A(_09595_),
    .B(_09600_),
    .Y(_09601_));
 sky130_fd_sc_hd__xor2_4 _26265_ (.A(_09594_),
    .B(_09601_),
    .X(_09602_));
 sky130_fd_sc_hd__xnor2_4 _26266_ (.A(_09593_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__xnor2_4 _26267_ (.A(_09591_),
    .B(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__and2_1 _26268_ (.A(_09394_),
    .B(_09392_),
    .X(_09605_));
 sky130_fd_sc_hd__o21ba_4 _26269_ (.A1(_09376_),
    .A2(_09395_),
    .B1_N(_09605_),
    .X(_09606_));
 sky130_fd_sc_hd__xor2_4 _26270_ (.A(_09604_),
    .B(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__xor2_4 _26271_ (.A(_09577_),
    .B(_09607_),
    .X(_09608_));
 sky130_fd_sc_hd__a21o_2 _26272_ (.A1(_09574_),
    .A2(_09575_),
    .B1(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__nand3_4 _26273_ (.A(_09574_),
    .B(_09608_),
    .C(_09575_),
    .Y(_09610_));
 sky130_fd_sc_hd__a21oi_2 _26274_ (.A1(_09398_),
    .A2(_09399_),
    .B1(_09400_),
    .Y(_09611_));
 sky130_fd_sc_hd__o21ai_4 _26275_ (.A1(_09437_),
    .A2(_09611_),
    .B1(_09402_),
    .Y(_09612_));
 sky130_fd_sc_hd__a21oi_4 _26276_ (.A1(_09609_),
    .A2(_09610_),
    .B1(_09612_),
    .Y(_09613_));
 sky130_fd_sc_hd__nand3_4 _26277_ (.A(_09612_),
    .B(_09609_),
    .C(_09610_),
    .Y(_09614_));
 sky130_vsdinv _26278_ (.A(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__and2_1 _26279_ (.A(_09461_),
    .B(_09452_),
    .X(_09616_));
 sky130_fd_sc_hd__nor2_1 _26280_ (.A(_09454_),
    .B(_09459_),
    .Y(_09617_));
 sky130_fd_sc_hd__o21ba_1 _26281_ (.A1(_09453_),
    .A2(_09460_),
    .B1_N(_09617_),
    .X(_09618_));
 sky130_fd_sc_hd__or2b_1 _26282_ (.A(_09417_),
    .B_N(_09409_),
    .X(_09619_));
 sky130_fd_sc_hd__o21ai_4 _26283_ (.A1(_09416_),
    .A2(_09410_),
    .B1(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__o21a_2 _26284_ (.A1(_09455_),
    .A2(_09458_),
    .B1(_09456_),
    .X(_09621_));
 sky130_fd_sc_hd__a2bb2oi_4 _26285_ (.A1_N(_14297_),
    .A2_N(_09406_),
    .B1(_09405_),
    .B2(_09407_),
    .Y(_09622_));
 sky130_fd_sc_hd__nand2_8 _26286_ (.A(_12776_),
    .B(_04996_),
    .Y(_09623_));
 sky130_fd_sc_hd__nand3_4 _26287_ (.A(_05131_),
    .B(_05064_),
    .C(_08077_),
    .Y(_09624_));
 sky130_fd_sc_hd__a22o_1 _26288_ (.A1(_05131_),
    .A2(_08077_),
    .B1(_05163_),
    .B2(_08170_),
    .X(_09625_));
 sky130_fd_sc_hd__o21ai_4 _26289_ (.A1(_14274_),
    .A2(_09624_),
    .B1(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__xnor2_4 _26290_ (.A(_09623_),
    .B(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__xnor2_4 _26291_ (.A(_09622_),
    .B(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__xor2_4 _26292_ (.A(_09621_),
    .B(_09628_),
    .X(_09629_));
 sky130_fd_sc_hd__xnor2_1 _26293_ (.A(_09620_),
    .B(_09629_),
    .Y(_09630_));
 sky130_fd_sc_hd__xor2_1 _26294_ (.A(_09618_),
    .B(_09630_),
    .X(_09631_));
 sky130_vsdinv _26295_ (.A(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__o21bai_1 _26296_ (.A1(_09616_),
    .A2(_09465_),
    .B1_N(_09632_),
    .Y(_09633_));
 sky130_vsdinv _26297_ (.A(_09616_),
    .Y(_09634_));
 sky130_fd_sc_hd__o211ai_2 _26298_ (.A1(_09450_),
    .A2(_09462_),
    .B1(_09634_),
    .C1(_09632_),
    .Y(_09635_));
 sky130_fd_sc_hd__o31ai_4 _26299_ (.A1(_05316_),
    .A2(_08604_),
    .A3(_04715_),
    .B1(_12781_),
    .Y(_09636_));
 sky130_fd_sc_hd__nor3_1 _26300_ (.A(_09636_),
    .B(_09472_),
    .C(_08987_),
    .Y(_09637_));
 sky130_fd_sc_hd__a21o_1 _26301_ (.A1(_08987_),
    .A2(_09636_),
    .B1(_09637_),
    .X(_09638_));
 sky130_fd_sc_hd__xor2_2 _26302_ (.A(_09278_),
    .B(_09638_),
    .X(_09639_));
 sky130_fd_sc_hd__a21o_1 _26303_ (.A1(_09633_),
    .A2(_09635_),
    .B1(_09639_),
    .X(_09640_));
 sky130_fd_sc_hd__and3_1 _26304_ (.A(_09633_),
    .B(_09639_),
    .C(_09635_),
    .X(_09641_));
 sky130_vsdinv _26305_ (.A(_09641_),
    .Y(_09642_));
 sky130_fd_sc_hd__or2b_1 _26306_ (.A(_09433_),
    .B_N(_09431_),
    .X(_09643_));
 sky130_fd_sc_hd__nand2_2 _26307_ (.A(_09435_),
    .B(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__a21o_1 _26308_ (.A1(_09640_),
    .A2(_09642_),
    .B1(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__nand3_4 _26309_ (.A(_09644_),
    .B(_09642_),
    .C(_09640_),
    .Y(_09646_));
 sky130_fd_sc_hd__a21boi_1 _26310_ (.A1(_09477_),
    .A2(_09467_),
    .B1_N(_09464_),
    .Y(_09647_));
 sky130_fd_sc_hd__a21bo_1 _26311_ (.A1(_09645_),
    .A2(_09646_),
    .B1_N(_09647_),
    .X(_09648_));
 sky130_fd_sc_hd__nand3b_4 _26312_ (.A_N(_09647_),
    .B(_09645_),
    .C(_09646_),
    .Y(_09649_));
 sky130_fd_sc_hd__nand2_4 _26313_ (.A(_09648_),
    .B(_09649_),
    .Y(_09650_));
 sky130_fd_sc_hd__o21ai_4 _26314_ (.A1(_09613_),
    .A2(_09615_),
    .B1(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__a21o_1 _26315_ (.A1(_09609_),
    .A2(_09610_),
    .B1(_09612_),
    .X(_09652_));
 sky130_fd_sc_hd__nand3b_4 _26316_ (.A_N(_09650_),
    .B(_09614_),
    .C(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__a21oi_4 _26317_ (.A1(_09444_),
    .A2(_09440_),
    .B1(_09442_),
    .Y(_09654_));
 sky130_fd_sc_hd__o21ai_4 _26318_ (.A1(_09489_),
    .A2(_09654_),
    .B1(_09445_),
    .Y(_09655_));
 sky130_fd_sc_hd__a21o_1 _26319_ (.A1(_09651_),
    .A2(_09653_),
    .B1(_09655_),
    .X(_09656_));
 sky130_fd_sc_hd__nand3_4 _26320_ (.A(_09655_),
    .B(_09651_),
    .C(_09653_),
    .Y(_09657_));
 sky130_fd_sc_hd__nand2_1 _26321_ (.A(_09475_),
    .B(_09473_),
    .Y(_09658_));
 sky130_fd_sc_hd__o21a_2 _26322_ (.A1(_09279_),
    .A2(_09476_),
    .B1(_09658_),
    .X(_09659_));
 sky130_fd_sc_hd__a21boi_4 _26323_ (.A1(_09482_),
    .A2(_09486_),
    .B1_N(_09483_),
    .Y(_09660_));
 sky130_fd_sc_hd__xor2_4 _26324_ (.A(_09659_),
    .B(_09660_),
    .X(_09661_));
 sky130_fd_sc_hd__a21oi_1 _26325_ (.A1(_09656_),
    .A2(_09657_),
    .B1(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__nand3_4 _26326_ (.A(_09656_),
    .B(_09661_),
    .C(_09657_),
    .Y(_09663_));
 sky130_vsdinv _26327_ (.A(_09663_),
    .Y(_09664_));
 sky130_vsdinv _26328_ (.A(_09498_),
    .Y(_09665_));
 sky130_fd_sc_hd__o21ai_4 _26329_ (.A1(_09665_),
    .A2(_09504_),
    .B1(_09494_),
    .Y(_09666_));
 sky130_fd_sc_hd__o21bai_2 _26330_ (.A1(_09662_),
    .A2(_09664_),
    .B1_N(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__a21oi_4 _26331_ (.A1(_09651_),
    .A2(_09653_),
    .B1(_09655_),
    .Y(_09668_));
 sky130_vsdinv _26332_ (.A(_09657_),
    .Y(_09669_));
 sky130_fd_sc_hd__o21bai_4 _26333_ (.A1(_09668_),
    .A2(_09669_),
    .B1_N(_09661_),
    .Y(_09670_));
 sky130_fd_sc_hd__nand3_4 _26334_ (.A(_09670_),
    .B(_09666_),
    .C(_09663_),
    .Y(_09671_));
 sky130_fd_sc_hd__a21boi_4 _26335_ (.A1(_09303_),
    .A2(_09299_),
    .B1_N(_09496_),
    .Y(_09672_));
 sky130_fd_sc_hd__a21oi_2 _26336_ (.A1(_09667_),
    .A2(_09671_),
    .B1(_09672_),
    .Y(_09673_));
 sky130_vsdinv _26337_ (.A(_09672_),
    .Y(_09674_));
 sky130_fd_sc_hd__a21oi_4 _26338_ (.A1(_09670_),
    .A2(_09663_),
    .B1(_09666_),
    .Y(_09675_));
 sky130_fd_sc_hd__nor3b_4 _26339_ (.A(_09674_),
    .B(_09675_),
    .C_N(_09671_),
    .Y(_09676_));
 sky130_fd_sc_hd__o21ai_2 _26340_ (.A1(_09509_),
    .A2(_09510_),
    .B1(_09507_),
    .Y(_09677_));
 sky130_fd_sc_hd__o21bai_4 _26341_ (.A1(_09673_),
    .A2(_09676_),
    .B1_N(_09677_),
    .Y(_09678_));
 sky130_fd_sc_hd__a21o_1 _26342_ (.A1(_09667_),
    .A2(_09671_),
    .B1(_09672_),
    .X(_09679_));
 sky130_fd_sc_hd__nand3_2 _26343_ (.A(_09667_),
    .B(_09672_),
    .C(_09671_),
    .Y(_09680_));
 sky130_fd_sc_hd__nand3_4 _26344_ (.A(_09679_),
    .B(_09677_),
    .C(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__nand2_4 _26345_ (.A(_09678_),
    .B(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__a21bo_1 _26346_ (.A1(_09335_),
    .A2(_09517_),
    .B1_N(_09513_),
    .X(_09683_));
 sky130_fd_sc_hd__o31ai_4 _26347_ (.A1(_09336_),
    .A2(_09518_),
    .A3(net409),
    .B1(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__xnor2_4 _26348_ (.A(_09682_),
    .B(_09684_),
    .Y(_02657_));
 sky130_fd_sc_hd__and2b_1 _26349_ (.A_N(_09545_),
    .B(_09528_),
    .X(_09685_));
 sky130_fd_sc_hd__o21a_2 _26350_ (.A1(_09522_),
    .A2(_09525_),
    .B1(_09523_),
    .X(_09686_));
 sky130_fd_sc_hd__a2bb2oi_4 _26351_ (.A1_N(_14401_),
    .A2_N(_09532_),
    .B1(_09531_),
    .B2(_09533_),
    .Y(_09687_));
 sky130_fd_sc_hd__nand2_2 _26352_ (.A(_07106_),
    .B(_05700_),
    .Y(_09688_));
 sky130_fd_sc_hd__or4_4 _26353_ (.A(_08402_),
    .B(_13989_),
    .C(_14377_),
    .D(_14382_),
    .X(_09689_));
 sky130_fd_sc_hd__a22o_1 _26354_ (.A1(_07262_),
    .A2(_06160_),
    .B1(_07102_),
    .B2(_09198_),
    .X(_09690_));
 sky130_fd_sc_hd__nand2_2 _26355_ (.A(_09689_),
    .B(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__xnor2_4 _26356_ (.A(_09688_),
    .B(_09691_),
    .Y(_09692_));
 sky130_fd_sc_hd__xnor2_4 _26357_ (.A(_09687_),
    .B(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__xor2_4 _26358_ (.A(_09686_),
    .B(_09693_),
    .X(_09694_));
 sky130_fd_sc_hd__or2b_1 _26359_ (.A(_09542_),
    .B_N(_09537_),
    .X(_09695_));
 sky130_fd_sc_hd__o21ai_4 _26360_ (.A1(_09535_),
    .A2(_09543_),
    .B1(_09695_),
    .Y(_09696_));
 sky130_fd_sc_hd__and2_2 _26361_ (.A(_07358_),
    .B(_05505_),
    .X(_09697_));
 sky130_fd_sc_hd__nand3_4 _26362_ (.A(_08374_),
    .B(_08375_),
    .C(_05405_),
    .Y(_09698_));
 sky130_fd_sc_hd__a22o_2 _26363_ (.A1(_07961_),
    .A2(_05405_),
    .B1(_08375_),
    .B2(_05497_),
    .X(_09699_));
 sky130_fd_sc_hd__o21ai_4 _26364_ (.A1(_05418_),
    .A2(_09698_),
    .B1(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__xor2_4 _26365_ (.A(_09697_),
    .B(_09700_),
    .X(_09701_));
 sky130_fd_sc_hd__nand3b_2 _26366_ (.A_N(_09539_),
    .B(_08526_),
    .C(_05057_),
    .Y(_09702_));
 sky130_fd_sc_hd__o31ai_4 _26367_ (.A1(_13966_),
    .A2(_14411_),
    .A3(_09541_),
    .B1(_09702_),
    .Y(_09703_));
 sky130_fd_sc_hd__and2_2 _26368_ (.A(_08644_),
    .B(_05308_),
    .X(_09704_));
 sky130_fd_sc_hd__nand2_2 _26369_ (.A(_08646_),
    .B(_05227_),
    .Y(_09705_));
 sky130_fd_sc_hd__and2b_2 _26370_ (.A_N(_05586_),
    .B(_08383_),
    .X(_09706_));
 sky130_fd_sc_hd__xor2_4 _26371_ (.A(_09705_),
    .B(_09706_),
    .X(_09707_));
 sky130_fd_sc_hd__xor2_4 _26372_ (.A(_09704_),
    .B(_09707_),
    .X(_09708_));
 sky130_fd_sc_hd__xor2_4 _26373_ (.A(_09703_),
    .B(_09708_),
    .X(_09709_));
 sky130_fd_sc_hd__xor2_4 _26374_ (.A(_09701_),
    .B(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__xnor2_2 _26375_ (.A(_09696_),
    .B(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__xnor2_2 _26376_ (.A(_09694_),
    .B(_09711_),
    .Y(_09712_));
 sky130_fd_sc_hd__a211o_2 _26377_ (.A1(_09544_),
    .A2(_09530_),
    .B1(_09685_),
    .C1(_09712_),
    .X(_09713_));
 sky130_fd_sc_hd__a21o_1 _26378_ (.A1(_09544_),
    .A2(_09530_),
    .B1(_09685_),
    .X(_09714_));
 sky130_fd_sc_hd__nand2_4 _26379_ (.A(_09714_),
    .B(_09712_),
    .Y(_09715_));
 sky130_fd_sc_hd__nor2_1 _26380_ (.A(_09521_),
    .B(_09526_),
    .Y(_09716_));
 sky130_fd_sc_hd__o21bai_2 _26381_ (.A1(_09520_),
    .A2(_09527_),
    .B1_N(_09716_),
    .Y(_09717_));
 sky130_fd_sc_hd__and2_2 _26382_ (.A(_08261_),
    .B(_06761_),
    .X(_09718_));
 sky130_fd_sc_hd__nand3_4 _26383_ (.A(_08422_),
    .B(_08859_),
    .C(_06584_),
    .Y(_09719_));
 sky130_fd_sc_hd__a22o_1 _26384_ (.A1(_08662_),
    .A2(_08342_),
    .B1(_09379_),
    .B2(_06441_),
    .X(_09720_));
 sky130_fd_sc_hd__o21ai_2 _26385_ (.A1(_14341_),
    .A2(_09719_),
    .B1(_09720_),
    .Y(_09721_));
 sky130_fd_sc_hd__xor2_2 _26386_ (.A(_09718_),
    .B(_09721_),
    .X(_09722_));
 sky130_fd_sc_hd__buf_4 _26387_ (.A(_07979_),
    .X(_09723_));
 sky130_fd_sc_hd__a22o_1 _26388_ (.A1(_07247_),
    .A2(_06019_),
    .B1(_09723_),
    .B2(_06030_),
    .X(_09724_));
 sky130_fd_sc_hd__nand3_4 _26389_ (.A(_08667_),
    .B(_08864_),
    .C(_05777_),
    .Y(_09725_));
 sky130_fd_sc_hd__or2b_1 _26390_ (.A(_09725_),
    .B_N(_06147_),
    .X(_09726_));
 sky130_fd_sc_hd__o2bb2ai_1 _26391_ (.A1_N(_09724_),
    .A2_N(_09726_),
    .B1(_14006_),
    .B2(_08338_),
    .Y(_09727_));
 sky130_fd_sc_hd__o2111ai_4 _26392_ (.A1(_06034_),
    .A2(_09725_),
    .B1(_09388_),
    .C1(_06280_),
    .D1(_09724_),
    .Y(_09728_));
 sky130_fd_sc_hd__nand2_2 _26393_ (.A(_09727_),
    .B(_09728_),
    .Y(_09729_));
 sky130_fd_sc_hd__o21a_1 _26394_ (.A1(_09562_),
    .A2(_09565_),
    .B1(_09563_),
    .X(_09730_));
 sky130_fd_sc_hd__xnor2_1 _26395_ (.A(_09729_),
    .B(_09730_),
    .Y(_09731_));
 sky130_fd_sc_hd__xor2_1 _26396_ (.A(_09722_),
    .B(_09731_),
    .X(_09732_));
 sky130_fd_sc_hd__or2_1 _26397_ (.A(_09717_),
    .B(_09732_),
    .X(_09733_));
 sky130_fd_sc_hd__nand2_1 _26398_ (.A(_09732_),
    .B(_09717_),
    .Y(_09734_));
 sky130_fd_sc_hd__nor2_1 _26399_ (.A(_09561_),
    .B(_09566_),
    .Y(_09735_));
 sky130_fd_sc_hd__o21bai_2 _26400_ (.A1(_09560_),
    .A2(_09567_),
    .B1_N(_09735_),
    .Y(_09736_));
 sky130_fd_sc_hd__a21oi_1 _26401_ (.A1(_09733_),
    .A2(_09734_),
    .B1(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__and3_1 _26402_ (.A(_09733_),
    .B(_09736_),
    .C(_09734_),
    .X(_09738_));
 sky130_fd_sc_hd__nor2_2 _26403_ (.A(_09737_),
    .B(_09738_),
    .Y(_09739_));
 sky130_fd_sc_hd__a21oi_1 _26404_ (.A1(_09713_),
    .A2(_09715_),
    .B1(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__nand3_4 _26405_ (.A(_09713_),
    .B(_09739_),
    .C(_09715_),
    .Y(_09741_));
 sky130_fd_sc_hd__nand2_2 _26406_ (.A(_09572_),
    .B(_09551_),
    .Y(_09742_));
 sky130_fd_sc_hd__nand3b_4 _26407_ (.A_N(_09740_),
    .B(_09741_),
    .C(_09742_),
    .Y(_09743_));
 sky130_vsdinv _26408_ (.A(_09740_),
    .Y(_09744_));
 sky130_fd_sc_hd__a21o_2 _26409_ (.A1(_09744_),
    .A2(_09741_),
    .B1(_09742_),
    .X(_09745_));
 sky130_fd_sc_hd__or2b_1 _26410_ (.A(_09603_),
    .B_N(_09591_),
    .X(_09746_));
 sky130_fd_sc_hd__nand2_1 _26411_ (.A(_09602_),
    .B(_09593_),
    .Y(_09747_));
 sky130_fd_sc_hd__and2_2 _26412_ (.A(_09746_),
    .B(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__o21a_2 _26413_ (.A1(_14309_),
    .A2(_09585_),
    .B1(_09588_),
    .X(_09749_));
 sky130_fd_sc_hd__a22o_1 _26414_ (.A1(_07281_),
    .A2(_07044_),
    .B1(_09071_),
    .B2(_07216_),
    .X(_09750_));
 sky130_fd_sc_hd__nand3_4 _26415_ (.A(_14037_),
    .B(_14042_),
    .C(_07209_),
    .Y(_09751_));
 sky130_fd_sc_hd__or2b_2 _26416_ (.A(_09751_),
    .B_N(_07477_),
    .X(_09752_));
 sky130_fd_sc_hd__o2bb2ai_1 _26417_ (.A1_N(_09750_),
    .A2_N(_09752_),
    .B1(_14048_),
    .B2(_14297_),
    .Y(_09753_));
 sky130_fd_sc_hd__o2111ai_4 _26418_ (.A1(_14303_),
    .A2(_09751_),
    .B1(_05442_),
    .C1(_07578_),
    .D1(_09750_),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2_2 _26419_ (.A(_09753_),
    .B(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__xnor2_4 _26420_ (.A(_09749_),
    .B(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__and2_2 _26421_ (.A(_05205_),
    .B(_08078_),
    .X(_09757_));
 sky130_fd_sc_hd__or4_4 _26422_ (.A(_14051_),
    .B(_14054_),
    .C(_14284_),
    .D(_14290_),
    .X(_09758_));
 sky130_fd_sc_hd__a22o_1 _26423_ (.A1(_05582_),
    .A2(_08779_),
    .B1(_05273_),
    .B2(_08487_),
    .X(_09759_));
 sky130_fd_sc_hd__nand2_2 _26424_ (.A(_09758_),
    .B(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__xor2_4 _26425_ (.A(_09757_),
    .B(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__xor2_4 _26426_ (.A(_09756_),
    .B(_09761_),
    .X(_09762_));
 sky130_fd_sc_hd__nor2_1 _26427_ (.A(_09595_),
    .B(_09600_),
    .Y(_09763_));
 sky130_fd_sc_hd__o21bai_4 _26428_ (.A1(_09594_),
    .A2(_09601_),
    .B1_N(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__a2bb2oi_4 _26429_ (.A1_N(_14329_),
    .A2_N(_09597_),
    .B1(_09596_),
    .B2(_09598_),
    .Y(_09765_));
 sky130_fd_sc_hd__a2bb2oi_4 _26430_ (.A1_N(_14347_),
    .A2_N(_09557_),
    .B1(_09556_),
    .B2(_09558_),
    .Y(_09766_));
 sky130_fd_sc_hd__and2_2 _26431_ (.A(_05717_),
    .B(_07039_),
    .X(_09767_));
 sky130_fd_sc_hd__nand3_4 _26432_ (.A(_05941_),
    .B(_05814_),
    .C(_06596_),
    .Y(_09768_));
 sky130_fd_sc_hd__a22o_2 _26433_ (.A1(_05943_),
    .A2(_06939_),
    .B1(_06071_),
    .B2(_07205_),
    .X(_09769_));
 sky130_fd_sc_hd__o21ai_4 _26434_ (.A1(_14320_),
    .A2(_09768_),
    .B1(_09769_),
    .Y(_09770_));
 sky130_fd_sc_hd__xor2_4 _26435_ (.A(_09767_),
    .B(_09770_),
    .X(_09771_));
 sky130_fd_sc_hd__xnor2_4 _26436_ (.A(_09766_),
    .B(_09771_),
    .Y(_09772_));
 sky130_fd_sc_hd__xor2_4 _26437_ (.A(_09765_),
    .B(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__xnor2_2 _26438_ (.A(_09764_),
    .B(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__xnor2_2 _26439_ (.A(_09762_),
    .B(_09774_),
    .Y(_09775_));
 sky130_fd_sc_hd__and2_1 _26440_ (.A(_09568_),
    .B(_09555_),
    .X(_09776_));
 sky130_fd_sc_hd__o21bai_4 _26441_ (.A1(_09553_),
    .A2(_09569_),
    .B1_N(_09776_),
    .Y(_09777_));
 sky130_fd_sc_hd__nor2_4 _26442_ (.A(_09775_),
    .B(_09777_),
    .Y(_09778_));
 sky130_fd_sc_hd__nand2_2 _26443_ (.A(_09777_),
    .B(_09775_),
    .Y(_09779_));
 sky130_fd_sc_hd__nor3b_4 _26444_ (.A(_09748_),
    .B(_09778_),
    .C_N(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__and2_1 _26445_ (.A(_09777_),
    .B(_09775_),
    .X(_09781_));
 sky130_fd_sc_hd__o21a_1 _26446_ (.A1(_09778_),
    .A2(_09781_),
    .B1(_09748_),
    .X(_09782_));
 sky130_fd_sc_hd__o2bb2ai_4 _26447_ (.A1_N(_09743_),
    .A2_N(_09745_),
    .B1(_09780_),
    .B2(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__nor2_2 _26448_ (.A(_09780_),
    .B(_09782_),
    .Y(_09784_));
 sky130_fd_sc_hd__nand3_4 _26449_ (.A(_09745_),
    .B(_09784_),
    .C(_09743_),
    .Y(_09785_));
 sky130_fd_sc_hd__nand2_2 _26450_ (.A(_09610_),
    .B(_09575_),
    .Y(_09786_));
 sky130_fd_sc_hd__a21o_1 _26451_ (.A1(_09783_),
    .A2(_09785_),
    .B1(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__nand3_4 _26452_ (.A(_09783_),
    .B(_09785_),
    .C(_09786_),
    .Y(_09788_));
 sky130_fd_sc_hd__or4_4 _26453_ (.A(_14075_),
    .B(_14098_),
    .C(_09284_),
    .D(_08987_),
    .X(_09789_));
 sky130_fd_sc_hd__o31ai_4 _26454_ (.A1(_08601_),
    .A2(_08986_),
    .A3(_09469_),
    .B1(_09789_),
    .Y(_09790_));
 sky130_fd_sc_hd__xor2_4 _26455_ (.A(_09278_),
    .B(_09790_),
    .X(_09791_));
 sky130_vsdinv _26456_ (.A(_09791_),
    .Y(_09792_));
 sky130_fd_sc_hd__buf_2 _26457_ (.A(_09792_),
    .X(_09793_));
 sky130_fd_sc_hd__nor2_2 _26458_ (.A(_09618_),
    .B(_09630_),
    .Y(_09794_));
 sky130_fd_sc_hd__a21oi_4 _26459_ (.A1(_09620_),
    .A2(_09629_),
    .B1(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__nor2_1 _26460_ (.A(_09622_),
    .B(_09627_),
    .Y(_09796_));
 sky130_fd_sc_hd__o21ba_2 _26461_ (.A1(_09621_),
    .A2(_09628_),
    .B1_N(_09796_),
    .X(_09797_));
 sky130_fd_sc_hd__or2b_1 _26462_ (.A(_09590_),
    .B_N(_09582_),
    .X(_09798_));
 sky130_fd_sc_hd__o21ai_4 _26463_ (.A1(_09589_),
    .A2(_09583_),
    .B1(_09798_),
    .Y(_09799_));
 sky130_fd_sc_hd__o22a_4 _26464_ (.A1(_14276_),
    .A2(_09624_),
    .B1(_09623_),
    .B2(_09626_),
    .X(_09800_));
 sky130_fd_sc_hd__a2bb2oi_4 _26465_ (.A1_N(_14291_),
    .A2_N(_09579_),
    .B1(_09578_),
    .B2(_09580_),
    .Y(_09801_));
 sky130_fd_sc_hd__nand2_2 _26466_ (.A(_14062_),
    .B(\pcpi_mul.rs1[31] ),
    .Y(_09802_));
 sky130_fd_sc_hd__nand2_8 _26467_ (.A(\pcpi_mul.rs1[32] ),
    .B(_05162_),
    .Y(_09803_));
 sky130_fd_sc_hd__xnor2_4 _26468_ (.A(_09802_),
    .B(_09803_),
    .Y(_09804_));
 sky130_fd_sc_hd__xnor2_4 _26469_ (.A(_09623_),
    .B(_09804_),
    .Y(_09805_));
 sky130_fd_sc_hd__xnor2_4 _26470_ (.A(_09801_),
    .B(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__xor2_4 _26471_ (.A(_09800_),
    .B(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__xnor2_4 _26472_ (.A(_09799_),
    .B(_09807_),
    .Y(_09808_));
 sky130_fd_sc_hd__xor2_4 _26473_ (.A(_09797_),
    .B(_09808_),
    .X(_09809_));
 sky130_fd_sc_hd__xor2_4 _26474_ (.A(_09795_),
    .B(_09809_),
    .X(_09810_));
 sky130_fd_sc_hd__nor2_2 _26475_ (.A(_09793_),
    .B(_09810_),
    .Y(_09811_));
 sky130_fd_sc_hd__and2_1 _26476_ (.A(_09810_),
    .B(_09793_),
    .X(_09812_));
 sky130_fd_sc_hd__or2b_2 _26477_ (.A(_09606_),
    .B_N(_09604_),
    .X(_09813_));
 sky130_fd_sc_hd__o221ai_4 _26478_ (.A1(_09577_),
    .A2(_09607_),
    .B1(_09811_),
    .B2(_09812_),
    .C1(_09813_),
    .Y(_09814_));
 sky130_fd_sc_hd__o21ai_1 _26479_ (.A1(_09577_),
    .A2(_09607_),
    .B1(_09813_),
    .Y(_09815_));
 sky130_vsdinv _26480_ (.A(_09811_),
    .Y(_09816_));
 sky130_fd_sc_hd__nand3b_2 _26481_ (.A_N(_09812_),
    .B(_09815_),
    .C(_09816_),
    .Y(_09817_));
 sky130_fd_sc_hd__a21boi_1 _26482_ (.A1(_09639_),
    .A2(_09635_),
    .B1_N(_09633_),
    .Y(_09818_));
 sky130_vsdinv _26483_ (.A(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__a21oi_2 _26484_ (.A1(_09814_),
    .A2(_09817_),
    .B1(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__and3_1 _26485_ (.A(_09814_),
    .B(_09817_),
    .C(_09819_),
    .X(_09821_));
 sky130_fd_sc_hd__nor2_4 _26486_ (.A(_09820_),
    .B(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__a21oi_1 _26487_ (.A1(_09787_),
    .A2(_09788_),
    .B1(_09822_),
    .Y(_09823_));
 sky130_vsdinv _26488_ (.A(_09822_),
    .Y(_09824_));
 sky130_fd_sc_hd__a21oi_4 _26489_ (.A1(_09783_),
    .A2(_09785_),
    .B1(_09786_),
    .Y(_09825_));
 sky130_fd_sc_hd__nor3b_4 _26490_ (.A(_09824_),
    .B(_09825_),
    .C_N(_09788_),
    .Y(_09826_));
 sky130_fd_sc_hd__o21ai_4 _26491_ (.A1(_09613_),
    .A2(_09650_),
    .B1(_09614_),
    .Y(_09827_));
 sky130_fd_sc_hd__o21bai_2 _26492_ (.A1(_09823_),
    .A2(_09826_),
    .B1_N(_09827_),
    .Y(_09828_));
 sky130_vsdinv _26493_ (.A(_09788_),
    .Y(_09829_));
 sky130_fd_sc_hd__o21bai_4 _26494_ (.A1(_09825_),
    .A2(_09829_),
    .B1_N(_09822_),
    .Y(_09830_));
 sky130_fd_sc_hd__nand3_4 _26495_ (.A(_09787_),
    .B(_09822_),
    .C(_09788_),
    .Y(_09831_));
 sky130_fd_sc_hd__nand3_4 _26496_ (.A(_09830_),
    .B(_09831_),
    .C(_09827_),
    .Y(_09832_));
 sky130_fd_sc_hd__o21ai_4 _26497_ (.A1(_09279_),
    .A2(_09638_),
    .B1(_09789_),
    .Y(_09833_));
 sky130_fd_sc_hd__nand2_2 _26498_ (.A(_09649_),
    .B(_09646_),
    .Y(_09834_));
 sky130_fd_sc_hd__xor2_4 _26499_ (.A(_09833_),
    .B(_09834_),
    .X(_09835_));
 sky130_fd_sc_hd__a21oi_1 _26500_ (.A1(_09828_),
    .A2(_09832_),
    .B1(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__nand3_4 _26501_ (.A(_09828_),
    .B(_09835_),
    .C(_09832_),
    .Y(_09837_));
 sky130_vsdinv _26502_ (.A(_09837_),
    .Y(_09838_));
 sky130_vsdinv _26503_ (.A(_09661_),
    .Y(_09839_));
 sky130_fd_sc_hd__o21ai_4 _26504_ (.A1(_09839_),
    .A2(_09668_),
    .B1(_09657_),
    .Y(_09840_));
 sky130_fd_sc_hd__o21bai_1 _26505_ (.A1(_09836_),
    .A2(_09838_),
    .B1_N(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__a21oi_4 _26506_ (.A1(_09830_),
    .A2(_09831_),
    .B1(_09827_),
    .Y(_09842_));
 sky130_vsdinv _26507_ (.A(_09832_),
    .Y(_09843_));
 sky130_fd_sc_hd__o21bai_4 _26508_ (.A1(_09842_),
    .A2(_09843_),
    .B1_N(_09835_),
    .Y(_09844_));
 sky130_fd_sc_hd__nand3_4 _26509_ (.A(_09844_),
    .B(_09837_),
    .C(_09840_),
    .Y(_09845_));
 sky130_fd_sc_hd__a21oi_4 _26510_ (.A1(_09488_),
    .A2(_09483_),
    .B1(_09659_),
    .Y(_09846_));
 sky130_fd_sc_hd__a21oi_1 _26511_ (.A1(_09841_),
    .A2(_09845_),
    .B1(_09846_),
    .Y(_09847_));
 sky130_vsdinv _26512_ (.A(_09846_),
    .Y(_09848_));
 sky130_fd_sc_hd__a21oi_4 _26513_ (.A1(_09844_),
    .A2(_09837_),
    .B1(_09840_),
    .Y(_09849_));
 sky130_vsdinv _26514_ (.A(_09845_),
    .Y(_09850_));
 sky130_fd_sc_hd__nor3_4 _26515_ (.A(_09848_),
    .B(_09849_),
    .C(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__o21ai_2 _26516_ (.A1(_09674_),
    .A2(_09675_),
    .B1(_09671_),
    .Y(_09852_));
 sky130_fd_sc_hd__o21bai_2 _26517_ (.A1(_09847_),
    .A2(_09851_),
    .B1_N(_09852_),
    .Y(_09853_));
 sky130_fd_sc_hd__o21bai_2 _26518_ (.A1(_09849_),
    .A2(_09850_),
    .B1_N(_09846_),
    .Y(_09854_));
 sky130_fd_sc_hd__nand3_2 _26519_ (.A(_09841_),
    .B(_09846_),
    .C(_09845_),
    .Y(_09855_));
 sky130_fd_sc_hd__nand3_4 _26520_ (.A(_09854_),
    .B(_09852_),
    .C(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__nand2_4 _26521_ (.A(_09853_),
    .B(_09856_),
    .Y(_09857_));
 sky130_vsdinv _26522_ (.A(_09681_),
    .Y(_09858_));
 sky130_fd_sc_hd__a21oi_4 _26523_ (.A1(_09684_),
    .A2(_09678_),
    .B1(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__xor2_4 _26524_ (.A(_09857_),
    .B(_09859_),
    .X(_02658_));
 sky130_fd_sc_hd__o21a_2 _26525_ (.A1(_09688_),
    .A2(_09691_),
    .B1(_09689_),
    .X(_09860_));
 sky130_fd_sc_hd__a2bb2oi_4 _26526_ (.A1_N(_14395_),
    .A2_N(_09698_),
    .B1(_09697_),
    .B2(_09699_),
    .Y(_09861_));
 sky130_fd_sc_hd__nand2_2 _26527_ (.A(_08400_),
    .B(_06020_),
    .Y(_09862_));
 sky130_fd_sc_hd__or4_4 _26528_ (.A(_08402_),
    .B(_13989_),
    .C(_14371_),
    .D(_06264_),
    .X(_09863_));
 sky130_fd_sc_hd__a22o_1 _26529_ (.A1(_07262_),
    .A2(_09198_),
    .B1(_08405_),
    .B2(_05769_),
    .X(_09864_));
 sky130_fd_sc_hd__nand2_2 _26530_ (.A(_09863_),
    .B(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__xnor2_4 _26531_ (.A(_09862_),
    .B(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__xnor2_4 _26532_ (.A(_09861_),
    .B(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__xnor2_4 _26533_ (.A(_09860_),
    .B(_09867_),
    .Y(_09868_));
 sky130_fd_sc_hd__or2b_1 _26534_ (.A(_09708_),
    .B_N(_09703_),
    .X(_09869_));
 sky130_fd_sc_hd__o21ai_4 _26535_ (.A1(_09701_),
    .A2(_09709_),
    .B1(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__and2_2 _26536_ (.A(_08634_),
    .B(_06161_),
    .X(_09871_));
 sky130_fd_sc_hd__nand3_4 _26537_ (.A(_08396_),
    .B(_13978_),
    .C(_05414_),
    .Y(_09872_));
 sky130_fd_sc_hd__a22o_2 _26538_ (.A1(_09357_),
    .A2(_05322_),
    .B1(_09162_),
    .B2(_05424_),
    .X(_09873_));
 sky130_fd_sc_hd__o21ai_4 _26539_ (.A1(_07668_),
    .A2(_09872_),
    .B1(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__xor2_4 _26540_ (.A(_09871_),
    .B(_09874_),
    .X(_09875_));
 sky130_fd_sc_hd__buf_6 _26541_ (.A(_09025_),
    .X(_09876_));
 sky130_fd_sc_hd__nand3b_2 _26542_ (.A_N(_09705_),
    .B(_09876_),
    .C(_14418_),
    .Y(_09877_));
 sky130_fd_sc_hd__o31ai_4 _26543_ (.A1(_13967_),
    .A2(_14406_),
    .A3(_09707_),
    .B1(_09877_),
    .Y(_09878_));
 sky130_fd_sc_hd__and2_2 _26544_ (.A(_09172_),
    .B(_05614_),
    .X(_09879_));
 sky130_fd_sc_hd__nand2_2 _26545_ (.A(_09174_),
    .B(_05181_),
    .Y(_09880_));
 sky130_fd_sc_hd__and2b_1 _26546_ (.A_N(_05105_),
    .B(_09176_),
    .X(_09881_));
 sky130_fd_sc_hd__xor2_4 _26547_ (.A(_09880_),
    .B(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__xor2_4 _26548_ (.A(_09879_),
    .B(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__xor2_4 _26549_ (.A(_09878_),
    .B(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__xor2_4 _26550_ (.A(_09875_),
    .B(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__xnor2_4 _26551_ (.A(_09870_),
    .B(_09885_),
    .Y(_09886_));
 sky130_fd_sc_hd__xor2_4 _26552_ (.A(_09868_),
    .B(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__and2b_1 _26553_ (.A_N(_09711_),
    .B(_09694_),
    .X(_09888_));
 sky130_fd_sc_hd__a21o_2 _26554_ (.A1(_09710_),
    .A2(_09696_),
    .B1(_09888_),
    .X(_09889_));
 sky130_fd_sc_hd__nor2_1 _26555_ (.A(_09887_),
    .B(_09889_),
    .Y(_09890_));
 sky130_vsdinv _26556_ (.A(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__nand2_4 _26557_ (.A(_09889_),
    .B(_09887_),
    .Y(_09892_));
 sky130_fd_sc_hd__nor2_1 _26558_ (.A(_09729_),
    .B(_09730_),
    .Y(_09893_));
 sky130_fd_sc_hd__o21ba_2 _26559_ (.A1(_09722_),
    .A2(_09731_),
    .B1_N(_09893_),
    .X(_09894_));
 sky130_fd_sc_hd__nor2_1 _26560_ (.A(_09687_),
    .B(_09692_),
    .Y(_09895_));
 sky130_fd_sc_hd__o21bai_4 _26561_ (.A1(_09686_),
    .A2(_09693_),
    .B1_N(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__and2_2 _26562_ (.A(_08261_),
    .B(_06940_),
    .X(_09897_));
 sky130_fd_sc_hd__nand3_4 _26563_ (.A(_08425_),
    .B(_08426_),
    .C(_07747_),
    .Y(_09898_));
 sky130_fd_sc_hd__a22o_2 _26564_ (.A1(_06895_),
    .A2(_06577_),
    .B1(_06896_),
    .B2(_06587_),
    .X(_09899_));
 sky130_fd_sc_hd__o21ai_4 _26565_ (.A1(_14334_),
    .A2(_09898_),
    .B1(_09899_),
    .Y(_09900_));
 sky130_fd_sc_hd__xor2_4 _26566_ (.A(_09897_),
    .B(_09900_),
    .X(_09901_));
 sky130_fd_sc_hd__o21a_2 _26567_ (.A1(_14360_),
    .A2(_09725_),
    .B1(_09728_),
    .X(_09902_));
 sky130_fd_sc_hd__nand2_2 _26568_ (.A(_08673_),
    .B(_06584_),
    .Y(_09903_));
 sky130_fd_sc_hd__or4_4 _26569_ (.A(_13999_),
    .B(_14002_),
    .C(_14351_),
    .D(_14358_),
    .X(_09904_));
 sky130_fd_sc_hd__a22o_1 _26570_ (.A1(_08431_),
    .A2(_07650_),
    .B1(_08864_),
    .B2(_06288_),
    .X(_09905_));
 sky130_fd_sc_hd__nand2_2 _26571_ (.A(_09904_),
    .B(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__xnor2_4 _26572_ (.A(_09903_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__xnor2_4 _26573_ (.A(_09902_),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__xor2_4 _26574_ (.A(_09901_),
    .B(_09908_),
    .X(_09909_));
 sky130_fd_sc_hd__xnor2_4 _26575_ (.A(_09896_),
    .B(_09909_),
    .Y(_09910_));
 sky130_fd_sc_hd__xor2_4 _26576_ (.A(_09894_),
    .B(_09910_),
    .X(_09911_));
 sky130_fd_sc_hd__a21oi_1 _26577_ (.A1(_09891_),
    .A2(_09892_),
    .B1(_09911_),
    .Y(_09912_));
 sky130_vsdinv _26578_ (.A(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__nand3b_4 _26579_ (.A_N(_09890_),
    .B(_09911_),
    .C(_09892_),
    .Y(_09914_));
 sky130_fd_sc_hd__nand2_4 _26580_ (.A(_09741_),
    .B(_09715_),
    .Y(_09915_));
 sky130_fd_sc_hd__a21o_1 _26581_ (.A1(_09913_),
    .A2(_09914_),
    .B1(_09915_),
    .X(_09916_));
 sky130_fd_sc_hd__nand3b_4 _26582_ (.A_N(_09912_),
    .B(_09914_),
    .C(_09915_),
    .Y(_09917_));
 sky130_fd_sc_hd__or2b_1 _26583_ (.A(_09774_),
    .B_N(_09762_),
    .X(_09918_));
 sky130_fd_sc_hd__nand2_1 _26584_ (.A(_09773_),
    .B(_09764_),
    .Y(_09919_));
 sky130_fd_sc_hd__and2_2 _26585_ (.A(_09918_),
    .B(_09919_),
    .X(_09920_));
 sky130_fd_sc_hd__nand2_2 _26586_ (.A(_09754_),
    .B(_09752_),
    .Y(_09921_));
 sky130_fd_sc_hd__and2_2 _26587_ (.A(_08710_),
    .B(_07585_),
    .X(_09922_));
 sky130_fd_sc_hd__nand3_4 _26588_ (.A(_14038_),
    .B(_14043_),
    .C(_07568_),
    .Y(_09923_));
 sky130_fd_sc_hd__a22o_2 _26589_ (.A1(_05956_),
    .A2(_07216_),
    .B1(_09071_),
    .B2(_07485_),
    .X(_09924_));
 sky130_fd_sc_hd__o21ai_4 _26590_ (.A1(_14297_),
    .A2(_09923_),
    .B1(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__xor2_4 _26591_ (.A(_09922_),
    .B(_09925_),
    .X(_09926_));
 sky130_fd_sc_hd__xor2_4 _26592_ (.A(_09921_),
    .B(_09926_),
    .X(_09927_));
 sky130_fd_sc_hd__and2_2 _26593_ (.A(_05720_),
    .B(_08171_),
    .X(_09928_));
 sky130_fd_sc_hd__or4_4 _26594_ (.A(_14051_),
    .B(_14054_),
    .C(_14278_),
    .D(_14285_),
    .X(_09929_));
 sky130_fd_sc_hd__a22o_1 _26595_ (.A1(_05362_),
    .A2(_08073_),
    .B1(_05364_),
    .B2(_08165_),
    .X(_09930_));
 sky130_fd_sc_hd__nand2_2 _26596_ (.A(_09929_),
    .B(_09930_),
    .Y(_09931_));
 sky130_fd_sc_hd__xor2_4 _26597_ (.A(_09928_),
    .B(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__xor2_4 _26598_ (.A(_09927_),
    .B(_09932_),
    .X(_09933_));
 sky130_fd_sc_hd__nor2_1 _26599_ (.A(_09766_),
    .B(_09771_),
    .Y(_09934_));
 sky130_fd_sc_hd__o21bai_4 _26600_ (.A1(_09765_),
    .A2(_09772_),
    .B1_N(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__a2bb2oi_4 _26601_ (.A1_N(_14322_),
    .A2_N(_09768_),
    .B1(_09767_),
    .B2(_09769_),
    .Y(_09936_));
 sky130_fd_sc_hd__a2bb2oi_4 _26602_ (.A1_N(_14341_),
    .A2_N(_09719_),
    .B1(_09718_),
    .B2(_09720_),
    .Y(_09937_));
 sky130_fd_sc_hd__and2_2 _26603_ (.A(_05717_),
    .B(_07210_),
    .X(_09938_));
 sky130_fd_sc_hd__nand3_4 _26604_ (.A(_05941_),
    .B(_05944_),
    .C(_07205_),
    .Y(_09939_));
 sky130_fd_sc_hd__a22o_2 _26605_ (.A1(_06067_),
    .A2(_06777_),
    .B1(_06071_),
    .B2(_06957_),
    .X(_09940_));
 sky130_fd_sc_hd__o21ai_4 _26606_ (.A1(_14314_),
    .A2(_09939_),
    .B1(_09940_),
    .Y(_09941_));
 sky130_fd_sc_hd__xor2_4 _26607_ (.A(_09938_),
    .B(_09941_),
    .X(_09942_));
 sky130_fd_sc_hd__xnor2_4 _26608_ (.A(_09937_),
    .B(_09942_),
    .Y(_09943_));
 sky130_fd_sc_hd__xor2_4 _26609_ (.A(_09936_),
    .B(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__xnor2_4 _26610_ (.A(_09935_),
    .B(_09944_),
    .Y(_09945_));
 sky130_fd_sc_hd__xnor2_4 _26611_ (.A(_09933_),
    .B(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__a21bo_2 _26612_ (.A1(_09733_),
    .A2(_09736_),
    .B1_N(_09734_),
    .X(_09947_));
 sky130_fd_sc_hd__xor2_4 _26613_ (.A(_09946_),
    .B(_09947_),
    .X(_09948_));
 sky130_fd_sc_hd__xor2_4 _26614_ (.A(_09920_),
    .B(_09948_),
    .X(_09949_));
 sky130_fd_sc_hd__a21boi_1 _26615_ (.A1(_09916_),
    .A2(_09917_),
    .B1_N(_09949_),
    .Y(_09950_));
 sky130_fd_sc_hd__a21oi_4 _26616_ (.A1(_09913_),
    .A2(_09914_),
    .B1(_09915_),
    .Y(_09951_));
 sky130_fd_sc_hd__nor3b_4 _26617_ (.A(_09949_),
    .B(_09951_),
    .C_N(_09917_),
    .Y(_09952_));
 sky130_fd_sc_hd__nand2_2 _26618_ (.A(_09785_),
    .B(_09743_),
    .Y(_09953_));
 sky130_fd_sc_hd__o21bai_2 _26619_ (.A1(_09950_),
    .A2(_09952_),
    .B1_N(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__nand2_1 _26620_ (.A(_09916_),
    .B(_09917_),
    .Y(_09955_));
 sky130_fd_sc_hd__nand2_2 _26621_ (.A(_09955_),
    .B(_09949_),
    .Y(_09956_));
 sky130_fd_sc_hd__nand3b_4 _26622_ (.A_N(_09949_),
    .B(_09916_),
    .C(_09917_),
    .Y(_09957_));
 sky130_fd_sc_hd__nand3_4 _26623_ (.A(_09956_),
    .B(_09957_),
    .C(_09953_),
    .Y(_09958_));
 sky130_fd_sc_hd__nor2_1 _26624_ (.A(_09801_),
    .B(_09805_),
    .Y(_09959_));
 sky130_fd_sc_hd__o21ba_1 _26625_ (.A1(_09800_),
    .A2(_09806_),
    .B1_N(_09959_),
    .X(_09960_));
 sky130_fd_sc_hd__nor2_1 _26626_ (.A(_09749_),
    .B(_09755_),
    .Y(_09961_));
 sky130_fd_sc_hd__o21bai_2 _26627_ (.A1(_09756_),
    .A2(_09761_),
    .B1_N(_09961_),
    .Y(_09962_));
 sky130_fd_sc_hd__nand3b_2 _26628_ (.A_N(_09803_),
    .B(_05337_),
    .C(_08596_),
    .Y(_09963_));
 sky130_fd_sc_hd__o21a_1 _26629_ (.A1(_09623_),
    .A2(_09804_),
    .B1(_09963_),
    .X(_09964_));
 sky130_fd_sc_hd__nand2_4 _26630_ (.A(\pcpi_mul.rs1[32] ),
    .B(_05588_),
    .Y(_09965_));
 sky130_fd_sc_hd__xnor2_4 _26631_ (.A(_09803_),
    .B(_09965_),
    .Y(_09966_));
 sky130_fd_sc_hd__xor2_4 _26632_ (.A(_09623_),
    .B(_09966_),
    .X(_09967_));
 sky130_fd_sc_hd__buf_6 _26633_ (.A(_09967_),
    .X(_09968_));
 sky130_fd_sc_hd__a21bo_1 _26634_ (.A1(_09759_),
    .A2(_09757_),
    .B1_N(_09758_),
    .X(_09969_));
 sky130_fd_sc_hd__xnor2_2 _26635_ (.A(_09968_),
    .B(_09969_),
    .Y(_09970_));
 sky130_fd_sc_hd__xor2_2 _26636_ (.A(_09964_),
    .B(_09970_),
    .X(_09971_));
 sky130_fd_sc_hd__xnor2_1 _26637_ (.A(_09962_),
    .B(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__xor2_1 _26638_ (.A(_09960_),
    .B(_09972_),
    .X(_09973_));
 sky130_fd_sc_hd__nor2_1 _26639_ (.A(_09797_),
    .B(_09808_),
    .Y(_09974_));
 sky130_fd_sc_hd__a21oi_2 _26640_ (.A1(_09799_),
    .A2(_09807_),
    .B1(_09974_),
    .Y(_09975_));
 sky130_fd_sc_hd__or2b_1 _26641_ (.A(_09973_),
    .B_N(_09975_),
    .X(_09976_));
 sky130_fd_sc_hd__or2b_1 _26642_ (.A(_09975_),
    .B_N(_09973_),
    .X(_09977_));
 sky130_fd_sc_hd__buf_6 _26643_ (.A(_09791_),
    .X(_09978_));
 sky130_fd_sc_hd__a21oi_2 _26644_ (.A1(_09976_),
    .A2(_09977_),
    .B1(_09978_),
    .Y(_09979_));
 sky130_fd_sc_hd__and3_1 _26645_ (.A(_09976_),
    .B(_09977_),
    .C(_09791_),
    .X(_09980_));
 sky130_vsdinv _26646_ (.A(_09980_),
    .Y(_09981_));
 sky130_fd_sc_hd__o21ai_4 _26647_ (.A1(_09748_),
    .A2(_09778_),
    .B1(_09779_),
    .Y(_09982_));
 sky130_fd_sc_hd__nand3b_4 _26648_ (.A_N(_09979_),
    .B(_09981_),
    .C(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__o21bai_2 _26649_ (.A1(_09979_),
    .A2(_09980_),
    .B1_N(_09982_),
    .Y(_09984_));
 sky130_fd_sc_hd__buf_2 _26650_ (.A(_09793_),
    .X(_09985_));
 sky130_fd_sc_hd__or2b_1 _26651_ (.A(_09795_),
    .B_N(_09809_),
    .X(_09986_));
 sky130_fd_sc_hd__o21a_1 _26652_ (.A1(_09985_),
    .A2(_09810_),
    .B1(_09986_),
    .X(_09987_));
 sky130_fd_sc_hd__a21bo_1 _26653_ (.A1(_09983_),
    .A2(_09984_),
    .B1_N(_09987_),
    .X(_09988_));
 sky130_fd_sc_hd__nand3b_4 _26654_ (.A_N(_09987_),
    .B(_09983_),
    .C(_09984_),
    .Y(_09989_));
 sky130_fd_sc_hd__nand2_2 _26655_ (.A(_09988_),
    .B(_09989_),
    .Y(_09990_));
 sky130_vsdinv _26656_ (.A(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__a21oi_1 _26657_ (.A1(_09954_),
    .A2(_09958_),
    .B1(_09991_),
    .Y(_09992_));
 sky130_fd_sc_hd__nand3_4 _26658_ (.A(_09954_),
    .B(_09991_),
    .C(_09958_),
    .Y(_09993_));
 sky130_vsdinv _26659_ (.A(_09993_),
    .Y(_09994_));
 sky130_fd_sc_hd__o21ai_4 _26660_ (.A1(_09824_),
    .A2(_09825_),
    .B1(_09788_),
    .Y(_09995_));
 sky130_fd_sc_hd__o21bai_2 _26661_ (.A1(_09992_),
    .A2(_09994_),
    .B1_N(_09995_),
    .Y(_09996_));
 sky130_fd_sc_hd__nand2_1 _26662_ (.A(_09954_),
    .B(_09958_),
    .Y(_09997_));
 sky130_fd_sc_hd__nand2_2 _26663_ (.A(_09997_),
    .B(_09990_),
    .Y(_09998_));
 sky130_fd_sc_hd__nand3_4 _26664_ (.A(_09998_),
    .B(_09993_),
    .C(_09995_),
    .Y(_09999_));
 sky130_fd_sc_hd__o21a_2 _26665_ (.A1(_09279_),
    .A2(_09790_),
    .B1(_09789_),
    .X(_10000_));
 sky130_vsdinv _26666_ (.A(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__a21bo_2 _26667_ (.A1(_09819_),
    .A2(_09814_),
    .B1_N(_09817_),
    .X(_10002_));
 sky130_fd_sc_hd__xor2_4 _26668_ (.A(_10001_),
    .B(_10002_),
    .X(_10003_));
 sky130_fd_sc_hd__a21oi_1 _26669_ (.A1(_09996_),
    .A2(_09999_),
    .B1(_10003_),
    .Y(_10004_));
 sky130_vsdinv _26670_ (.A(_10003_),
    .Y(_10005_));
 sky130_fd_sc_hd__a21oi_4 _26671_ (.A1(_09998_),
    .A2(_09993_),
    .B1(_09995_),
    .Y(_10006_));
 sky130_fd_sc_hd__nor3b_2 _26672_ (.A(_10005_),
    .B(_10006_),
    .C_N(_09999_),
    .Y(_10007_));
 sky130_vsdinv _26673_ (.A(_09835_),
    .Y(_10008_));
 sky130_fd_sc_hd__o21ai_4 _26674_ (.A1(_10008_),
    .A2(_09842_),
    .B1(_09832_),
    .Y(_10009_));
 sky130_fd_sc_hd__o21bai_1 _26675_ (.A1(_10004_),
    .A2(_10007_),
    .B1_N(_10009_),
    .Y(_10010_));
 sky130_fd_sc_hd__and3_1 _26676_ (.A(_09998_),
    .B(_09993_),
    .C(_09995_),
    .X(_10011_));
 sky130_fd_sc_hd__o21bai_4 _26677_ (.A1(_10006_),
    .A2(_10011_),
    .B1_N(_10003_),
    .Y(_10012_));
 sky130_fd_sc_hd__nand3_4 _26678_ (.A(_09996_),
    .B(_10003_),
    .C(_09999_),
    .Y(_10013_));
 sky130_fd_sc_hd__nand3_4 _26679_ (.A(_10012_),
    .B(_10013_),
    .C(_10009_),
    .Y(_10014_));
 sky130_fd_sc_hd__a21boi_4 _26680_ (.A1(_09649_),
    .A2(_09646_),
    .B1_N(_09833_),
    .Y(_10015_));
 sky130_fd_sc_hd__a21oi_1 _26681_ (.A1(_10010_),
    .A2(_10014_),
    .B1(_10015_),
    .Y(_10016_));
 sky130_vsdinv _26682_ (.A(_10015_),
    .Y(_10017_));
 sky130_fd_sc_hd__a21oi_4 _26683_ (.A1(_10012_),
    .A2(_10013_),
    .B1(_10009_),
    .Y(_10018_));
 sky130_vsdinv _26684_ (.A(_10014_),
    .Y(_10019_));
 sky130_fd_sc_hd__nor3_1 _26685_ (.A(_10017_),
    .B(_10018_),
    .C(_10019_),
    .Y(_10020_));
 sky130_fd_sc_hd__o21ai_2 _26686_ (.A1(_09848_),
    .A2(_09849_),
    .B1(_09845_),
    .Y(_10021_));
 sky130_fd_sc_hd__o21bai_1 _26687_ (.A1(_10016_),
    .A2(_10020_),
    .B1_N(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__o21bai_2 _26688_ (.A1(_10018_),
    .A2(_10019_),
    .B1_N(_10015_),
    .Y(_10023_));
 sky130_fd_sc_hd__nand3_2 _26689_ (.A(_10010_),
    .B(_10015_),
    .C(_10014_),
    .Y(_10024_));
 sky130_fd_sc_hd__nand3_4 _26690_ (.A(_10023_),
    .B(_10024_),
    .C(_10021_),
    .Y(_10025_));
 sky130_fd_sc_hd__nand2_2 _26691_ (.A(_10022_),
    .B(_10025_),
    .Y(_10026_));
 sky130_fd_sc_hd__nor2_2 _26692_ (.A(_09336_),
    .B(_09518_),
    .Y(_10027_));
 sky130_fd_sc_hd__nor2_4 _26693_ (.A(_09682_),
    .B(_09857_),
    .Y(_10028_));
 sky130_fd_sc_hd__nand2_4 _26694_ (.A(_10027_),
    .B(_10028_),
    .Y(_10029_));
 sky130_fd_sc_hd__nor2_8 _26695_ (.A(_10029_),
    .B(_09340_),
    .Y(_10030_));
 sky130_fd_sc_hd__nor2_2 _26696_ (.A(_09145_),
    .B(_09146_),
    .Y(_10031_));
 sky130_fd_sc_hd__a31oi_4 _26697_ (.A1(_09144_),
    .A2(_10031_),
    .A3(_08959_),
    .B1(_09339_),
    .Y(_10032_));
 sky130_fd_sc_hd__a21boi_1 _26698_ (.A1(_09335_),
    .A2(_09517_),
    .B1_N(_09513_),
    .Y(_10033_));
 sky130_fd_sc_hd__a21bo_1 _26699_ (.A1(_09858_),
    .A2(_09853_),
    .B1_N(_09856_),
    .X(_10034_));
 sky130_fd_sc_hd__a21oi_2 _26700_ (.A1(_10028_),
    .A2(_10033_),
    .B1(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__o21ai_4 _26701_ (.A1(_10029_),
    .A2(_10032_),
    .B1(_10035_),
    .Y(_10036_));
 sky130_fd_sc_hd__a21oi_4 _26702_ (.A1(_08567_),
    .A2(_10030_),
    .B1(_10036_),
    .Y(_10037_));
 sky130_fd_sc_hd__xor2_1 _26703_ (.A(_10026_),
    .B(_10037_),
    .X(_02659_));
 sky130_fd_sc_hd__nor2_1 _26704_ (.A(_09902_),
    .B(_09907_),
    .Y(_10038_));
 sky130_fd_sc_hd__o21ba_1 _26705_ (.A1(_09901_),
    .A2(_09908_),
    .B1_N(_10038_),
    .X(_10039_));
 sky130_fd_sc_hd__nor2_1 _26706_ (.A(_09861_),
    .B(_09866_),
    .Y(_10040_));
 sky130_fd_sc_hd__o21bai_4 _26707_ (.A1(_09860_),
    .A2(_09867_),
    .B1_N(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__and2_2 _26708_ (.A(_06059_),
    .B(_07205_),
    .X(_10042_));
 sky130_fd_sc_hd__nand3_4 _26709_ (.A(_08662_),
    .B(_06896_),
    .C(_06450_),
    .Y(_10043_));
 sky130_fd_sc_hd__a22o_2 _26710_ (.A1(_14010_),
    .A2(_06587_),
    .B1(_14015_),
    .B2(_07033_),
    .X(_10044_));
 sky130_fd_sc_hd__o21ai_4 _26711_ (.A1(_14328_),
    .A2(_10043_),
    .B1(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__xor2_4 _26712_ (.A(_10042_),
    .B(_10045_),
    .X(_10046_));
 sky130_fd_sc_hd__and2_2 _26713_ (.A(_06649_),
    .B(_06577_),
    .X(_10047_));
 sky130_fd_sc_hd__nand3_4 _26714_ (.A(_08667_),
    .B(_08432_),
    .C(_06288_),
    .Y(_10048_));
 sky130_fd_sc_hd__a22o_2 _26715_ (.A1(_07246_),
    .A2(_06037_),
    .B1(_06647_),
    .B2(_06583_),
    .X(_10049_));
 sky130_fd_sc_hd__o21ai_4 _26716_ (.A1(_06293_),
    .A2(_10048_),
    .B1(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__xor2_4 _26717_ (.A(_10047_),
    .B(_10050_),
    .X(_10051_));
 sky130_fd_sc_hd__o21a_2 _26718_ (.A1(_09903_),
    .A2(_09906_),
    .B1(_09904_),
    .X(_10052_));
 sky130_fd_sc_hd__xnor2_4 _26719_ (.A(_10051_),
    .B(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__xor2_4 _26720_ (.A(_10046_),
    .B(_10053_),
    .X(_10054_));
 sky130_fd_sc_hd__xnor2_2 _26721_ (.A(_10041_),
    .B(_10054_),
    .Y(_10055_));
 sky130_fd_sc_hd__xor2_1 _26722_ (.A(_10039_),
    .B(_10055_),
    .X(_10056_));
 sky130_vsdinv _26723_ (.A(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__and2_1 _26724_ (.A(_09885_),
    .B(_09870_),
    .X(_10058_));
 sky130_fd_sc_hd__o21bai_4 _26725_ (.A1(_09868_),
    .A2(_09886_),
    .B1_N(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__o21a_2 _26726_ (.A1(_09862_),
    .A2(_09865_),
    .B1(_09863_),
    .X(_10060_));
 sky130_fd_sc_hd__a2bb2oi_4 _26727_ (.A1_N(_14390_),
    .A2_N(_09872_),
    .B1(_09871_),
    .B2(_09873_),
    .Y(_10061_));
 sky130_fd_sc_hd__and2_2 _26728_ (.A(_06887_),
    .B(_06030_),
    .X(_10062_));
 sky130_fd_sc_hd__nand3_4 _26729_ (.A(_08404_),
    .B(_08405_),
    .C(_05769_),
    .Y(_10063_));
 sky130_fd_sc_hd__a22o_2 _26730_ (.A1(_07262_),
    .A2(_05699_),
    .B1(_07102_),
    .B2(_05777_),
    .X(_10064_));
 sky130_fd_sc_hd__o21ai_4 _26731_ (.A1(_14366_),
    .A2(_10063_),
    .B1(_10064_),
    .Y(_10065_));
 sky130_fd_sc_hd__xor2_4 _26732_ (.A(_10062_),
    .B(_10065_),
    .X(_10066_));
 sky130_fd_sc_hd__xnor2_4 _26733_ (.A(_10061_),
    .B(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__xnor2_4 _26734_ (.A(_10060_),
    .B(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__or2b_1 _26735_ (.A(_09883_),
    .B_N(_09878_),
    .X(_10069_));
 sky130_fd_sc_hd__o21ai_4 _26736_ (.A1(_09875_),
    .A2(_09884_),
    .B1(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__and2_2 _26737_ (.A(_08634_),
    .B(_05611_),
    .X(_10071_));
 sky130_fd_sc_hd__nand3_4 _26738_ (.A(_09357_),
    .B(_08637_),
    .C(_05424_),
    .Y(_10072_));
 sky130_fd_sc_hd__a22o_2 _26739_ (.A1(_08374_),
    .A2(_05424_),
    .B1(_09164_),
    .B2(_05513_),
    .X(_10073_));
 sky130_fd_sc_hd__o21ai_4 _26740_ (.A1(_06409_),
    .A2(_10072_),
    .B1(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__xor2_4 _26741_ (.A(_10071_),
    .B(_10074_),
    .X(_10075_));
 sky130_fd_sc_hd__nand3b_2 _26742_ (.A_N(_09880_),
    .B(_08526_),
    .C(_14411_),
    .Y(_10076_));
 sky130_fd_sc_hd__o31ai_4 _26743_ (.A1(_09168_),
    .A2(_05874_),
    .A3(_09882_),
    .B1(_10076_),
    .Y(_10077_));
 sky130_fd_sc_hd__and2_2 _26744_ (.A(_08644_),
    .B(_05413_),
    .X(_10078_));
 sky130_fd_sc_hd__nand2_2 _26745_ (.A(_09174_),
    .B(_05613_),
    .Y(_10079_));
 sky130_fd_sc_hd__and2b_1 _26746_ (.A_N(_05236_),
    .B(_09176_),
    .X(_10080_));
 sky130_fd_sc_hd__xor2_4 _26747_ (.A(_10079_),
    .B(_10080_),
    .X(_10081_));
 sky130_fd_sc_hd__xor2_4 _26748_ (.A(_10078_),
    .B(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__xor2_4 _26749_ (.A(_10077_),
    .B(_10082_),
    .X(_10083_));
 sky130_fd_sc_hd__xor2_4 _26750_ (.A(_10075_),
    .B(_10083_),
    .X(_10084_));
 sky130_fd_sc_hd__xnor2_4 _26751_ (.A(_10070_),
    .B(_10084_),
    .Y(_10085_));
 sky130_fd_sc_hd__xor2_4 _26752_ (.A(_10068_),
    .B(_10085_),
    .X(_10086_));
 sky130_fd_sc_hd__xnor2_4 _26753_ (.A(_10059_),
    .B(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__nor2_2 _26754_ (.A(_10057_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__and2_1 _26755_ (.A(_10087_),
    .B(_10057_),
    .X(_10089_));
 sky130_fd_sc_hd__o211ai_4 _26756_ (.A1(_10088_),
    .A2(_10089_),
    .B1(_09892_),
    .C1(_09914_),
    .Y(_10090_));
 sky130_vsdinv _26757_ (.A(_10088_),
    .Y(_10091_));
 sky130_fd_sc_hd__nand2_1 _26758_ (.A(_09914_),
    .B(_09892_),
    .Y(_10092_));
 sky130_fd_sc_hd__nand3b_4 _26759_ (.A_N(_10089_),
    .B(_10091_),
    .C(_10092_),
    .Y(_10093_));
 sky130_fd_sc_hd__or2b_1 _26760_ (.A(_09945_),
    .B_N(_09933_),
    .X(_10094_));
 sky130_fd_sc_hd__a21boi_4 _26761_ (.A1(_09944_),
    .A2(_09935_),
    .B1_N(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__a2bb2oi_4 _26762_ (.A1_N(_14298_),
    .A2_N(_09923_),
    .B1(_09922_),
    .B2(_09924_),
    .Y(_10096_));
 sky130_fd_sc_hd__and2_2 _26763_ (.A(_08710_),
    .B(_08487_),
    .X(_10097_));
 sky130_fd_sc_hd__nand3_4 _26764_ (.A(_05956_),
    .B(_09071_),
    .C(_08782_),
    .Y(_10098_));
 sky130_fd_sc_hd__a22o_2 _26765_ (.A1(_07655_),
    .A2(_07484_),
    .B1(_05531_),
    .B2(_07584_),
    .X(_10099_));
 sky130_fd_sc_hd__o21ai_4 _26766_ (.A1(_14291_),
    .A2(_10098_),
    .B1(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__xor2_4 _26767_ (.A(_10097_),
    .B(_10100_),
    .X(_10101_));
 sky130_fd_sc_hd__xnor2_4 _26768_ (.A(_10096_),
    .B(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__and2_1 _26769_ (.A(\pcpi_mul.rs1[32] ),
    .B(\pcpi_mul.rs2[9] ),
    .X(_10103_));
 sky130_fd_sc_hd__buf_4 _26770_ (.A(_10103_),
    .X(_10104_));
 sky130_fd_sc_hd__or4_4 _26771_ (.A(_14051_),
    .B(_14054_),
    .C(_14274_),
    .D(_14278_),
    .X(_10105_));
 sky130_fd_sc_hd__a22o_1 _26772_ (.A1(_05581_),
    .A2(_08078_),
    .B1(_06200_),
    .B2(_08170_),
    .X(_10106_));
 sky130_fd_sc_hd__nand2_4 _26773_ (.A(_10105_),
    .B(_10106_),
    .Y(_10107_));
 sky130_fd_sc_hd__xor2_4 _26774_ (.A(_10104_),
    .B(_10107_),
    .X(_10108_));
 sky130_fd_sc_hd__xor2_4 _26775_ (.A(_10102_),
    .B(_10108_),
    .X(_10109_));
 sky130_fd_sc_hd__nor2_1 _26776_ (.A(_09937_),
    .B(_09942_),
    .Y(_10110_));
 sky130_fd_sc_hd__o21bai_4 _26777_ (.A1(_09936_),
    .A2(_09943_),
    .B1_N(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__a2bb2oi_4 _26778_ (.A1_N(_08464_),
    .A2_N(_09939_),
    .B1(_09938_),
    .B2(_09940_),
    .Y(_10112_));
 sky130_fd_sc_hd__a2bb2oi_4 _26779_ (.A1_N(_14334_),
    .A2_N(_09898_),
    .B1(_09897_),
    .B2(_09899_),
    .Y(_10113_));
 sky130_fd_sc_hd__and2_2 _26780_ (.A(_06355_),
    .B(_07568_),
    .X(_10114_));
 sky130_fd_sc_hd__nand3_4 _26781_ (.A(_06067_),
    .B(_08355_),
    .C(_06957_),
    .Y(_10115_));
 sky130_fd_sc_hd__a22o_2 _26782_ (.A1(_08354_),
    .A2(_07038_),
    .B1(_08357_),
    .B2(_07209_),
    .X(_10116_));
 sky130_fd_sc_hd__o21ai_4 _26783_ (.A1(_14308_),
    .A2(_10115_),
    .B1(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__xor2_4 _26784_ (.A(_10114_),
    .B(_10117_),
    .X(_10118_));
 sky130_fd_sc_hd__xnor2_4 _26785_ (.A(_10113_),
    .B(_10118_),
    .Y(_10119_));
 sky130_fd_sc_hd__xor2_4 _26786_ (.A(_10112_),
    .B(_10119_),
    .X(_10120_));
 sky130_fd_sc_hd__xnor2_4 _26787_ (.A(_10111_),
    .B(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__xnor2_4 _26788_ (.A(_10109_),
    .B(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__and2_1 _26789_ (.A(_09909_),
    .B(_09896_),
    .X(_10123_));
 sky130_fd_sc_hd__o21ba_4 _26790_ (.A1(_09894_),
    .A2(_09910_),
    .B1_N(_10123_),
    .X(_10124_));
 sky130_fd_sc_hd__xor2_4 _26791_ (.A(_10122_),
    .B(_10124_),
    .X(_10125_));
 sky130_fd_sc_hd__xor2_4 _26792_ (.A(_10095_),
    .B(_10125_),
    .X(_10126_));
 sky130_fd_sc_hd__a21oi_2 _26793_ (.A1(_10090_),
    .A2(_10093_),
    .B1(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__nand3_4 _26794_ (.A(_10126_),
    .B(_10090_),
    .C(_10093_),
    .Y(_10128_));
 sky130_vsdinv _26795_ (.A(_10128_),
    .Y(_10129_));
 sky130_fd_sc_hd__o21ai_2 _26796_ (.A1(_09949_),
    .A2(_09951_),
    .B1(_09917_),
    .Y(_10130_));
 sky130_fd_sc_hd__o21bai_2 _26797_ (.A1(_10127_),
    .A2(_10129_),
    .B1_N(_10130_),
    .Y(_10131_));
 sky130_fd_sc_hd__nand3b_4 _26798_ (.A_N(_10127_),
    .B(_10130_),
    .C(_10128_),
    .Y(_10132_));
 sky130_fd_sc_hd__nand2_1 _26799_ (.A(_09971_),
    .B(_09962_),
    .Y(_10133_));
 sky130_fd_sc_hd__o21a_1 _26800_ (.A1(_09960_),
    .A2(_09972_),
    .B1(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__buf_2 _26801_ (.A(_09968_),
    .X(_10135_));
 sky130_fd_sc_hd__nand2_1 _26802_ (.A(_09969_),
    .B(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__o21a_2 _26803_ (.A1(_09964_),
    .A2(_09970_),
    .B1(_10136_),
    .X(_10137_));
 sky130_fd_sc_hd__a21oi_1 _26804_ (.A1(_09752_),
    .A2(_09754_),
    .B1(_09926_),
    .Y(_10138_));
 sky130_fd_sc_hd__o21bai_4 _26805_ (.A1(_09927_),
    .A2(_09932_),
    .B1_N(_10138_),
    .Y(_10139_));
 sky130_fd_sc_hd__nand3_2 _26806_ (.A(_12778_),
    .B(_05127_),
    .C(_05065_),
    .Y(_10140_));
 sky130_fd_sc_hd__o21a_2 _26807_ (.A1(_09623_),
    .A2(_09966_),
    .B1(_10140_),
    .X(_10141_));
 sky130_fd_sc_hd__buf_6 _26808_ (.A(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__a21bo_2 _26809_ (.A1(_09930_),
    .A2(_09928_),
    .B1_N(_09929_),
    .X(_10143_));
 sky130_fd_sc_hd__xnor2_4 _26810_ (.A(_09968_),
    .B(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__xor2_4 _26811_ (.A(_10142_),
    .B(_10144_),
    .X(_10145_));
 sky130_fd_sc_hd__xnor2_4 _26812_ (.A(_10139_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__xor2_4 _26813_ (.A(_10137_),
    .B(_10146_),
    .X(_10147_));
 sky130_fd_sc_hd__xor2_2 _26814_ (.A(_10134_),
    .B(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__clkbuf_2 _26815_ (.A(_09792_),
    .X(_10149_));
 sky130_fd_sc_hd__and2_1 _26816_ (.A(_10148_),
    .B(_10149_),
    .X(_10150_));
 sky130_vsdinv _26817_ (.A(_09920_),
    .Y(_10151_));
 sky130_fd_sc_hd__and2_1 _26818_ (.A(_09947_),
    .B(_09946_),
    .X(_10152_));
 sky130_fd_sc_hd__a21o_1 _26819_ (.A1(_09948_),
    .A2(_10151_),
    .B1(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__nor2_1 _26820_ (.A(_09985_),
    .B(_10148_),
    .Y(_10154_));
 sky130_vsdinv _26821_ (.A(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__nand3b_4 _26822_ (.A_N(_10150_),
    .B(_10153_),
    .C(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__o21bai_2 _26823_ (.A1(_10154_),
    .A2(_10150_),
    .B1_N(_10153_),
    .Y(_10157_));
 sky130_fd_sc_hd__a21boi_1 _26824_ (.A1(_09978_),
    .A2(_09976_),
    .B1_N(_09977_),
    .Y(_10158_));
 sky130_fd_sc_hd__a21bo_1 _26825_ (.A1(_10156_),
    .A2(_10157_),
    .B1_N(_10158_),
    .X(_10159_));
 sky130_fd_sc_hd__nand3b_4 _26826_ (.A_N(_10158_),
    .B(_10156_),
    .C(_10157_),
    .Y(_10160_));
 sky130_fd_sc_hd__nand2_2 _26827_ (.A(_10159_),
    .B(_10160_),
    .Y(_10161_));
 sky130_vsdinv _26828_ (.A(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__a21o_1 _26829_ (.A1(_10131_),
    .A2(_10132_),
    .B1(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__nand3b_4 _26830_ (.A_N(_10161_),
    .B(_10131_),
    .C(_10132_),
    .Y(_10164_));
 sky130_fd_sc_hd__a21oi_2 _26831_ (.A1(_09956_),
    .A2(_09957_),
    .B1(_09953_),
    .Y(_10165_));
 sky130_fd_sc_hd__o21ai_4 _26832_ (.A1(_09990_),
    .A2(_10165_),
    .B1(_09958_),
    .Y(_10166_));
 sky130_fd_sc_hd__a21oi_4 _26833_ (.A1(_10163_),
    .A2(_10164_),
    .B1(_10166_),
    .Y(_10167_));
 sky130_fd_sc_hd__nand3_4 _26834_ (.A(_10163_),
    .B(_10166_),
    .C(_10164_),
    .Y(_10168_));
 sky130_vsdinv _26835_ (.A(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__buf_2 _26836_ (.A(_10001_),
    .X(_10170_));
 sky130_fd_sc_hd__nand2_2 _26837_ (.A(_09989_),
    .B(_09983_),
    .Y(_10171_));
 sky130_fd_sc_hd__xor2_4 _26838_ (.A(_10170_),
    .B(_10171_),
    .X(_10172_));
 sky130_fd_sc_hd__o21bai_4 _26839_ (.A1(_10167_),
    .A2(_10169_),
    .B1_N(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__nand3b_4 _26840_ (.A_N(_10167_),
    .B(_10172_),
    .C(_10168_),
    .Y(_10174_));
 sky130_fd_sc_hd__o21ai_4 _26841_ (.A1(_10005_),
    .A2(_10006_),
    .B1(_09999_),
    .Y(_10175_));
 sky130_fd_sc_hd__a21o_1 _26842_ (.A1(_10173_),
    .A2(_10174_),
    .B1(_10175_),
    .X(_10176_));
 sky130_fd_sc_hd__nand3_4 _26843_ (.A(_10173_),
    .B(_10174_),
    .C(_10175_),
    .Y(_10177_));
 sky130_fd_sc_hd__buf_6 _26844_ (.A(net414),
    .X(_10178_));
 sky130_fd_sc_hd__and2_1 _26845_ (.A(_10002_),
    .B(_10178_),
    .X(_10179_));
 sky130_fd_sc_hd__a21oi_1 _26846_ (.A1(_10176_),
    .A2(_10177_),
    .B1(_10179_),
    .Y(_10180_));
 sky130_vsdinv _26847_ (.A(_10179_),
    .Y(_10181_));
 sky130_fd_sc_hd__a21oi_4 _26848_ (.A1(_10173_),
    .A2(_10174_),
    .B1(_10175_),
    .Y(_10182_));
 sky130_vsdinv _26849_ (.A(_10177_),
    .Y(_10183_));
 sky130_fd_sc_hd__nor3_2 _26850_ (.A(_10181_),
    .B(_10182_),
    .C(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__o21ai_2 _26851_ (.A1(_10017_),
    .A2(_10018_),
    .B1(_10014_),
    .Y(_10185_));
 sky130_fd_sc_hd__o21bai_1 _26852_ (.A1(_10180_),
    .A2(_10184_),
    .B1_N(_10185_),
    .Y(_10186_));
 sky130_fd_sc_hd__o21bai_1 _26853_ (.A1(_10182_),
    .A2(_10183_),
    .B1_N(_10179_),
    .Y(_10187_));
 sky130_fd_sc_hd__nand3_2 _26854_ (.A(_10176_),
    .B(_10179_),
    .C(_10177_),
    .Y(_10188_));
 sky130_fd_sc_hd__nand3_2 _26855_ (.A(_10187_),
    .B(_10185_),
    .C(_10188_),
    .Y(_10189_));
 sky130_fd_sc_hd__nand2_2 _26856_ (.A(_10186_),
    .B(_10189_),
    .Y(_10190_));
 sky130_fd_sc_hd__o21a_1 _26857_ (.A1(_10026_),
    .A2(_10037_),
    .B1(_10025_),
    .X(_10191_));
 sky130_fd_sc_hd__xor2_1 _26858_ (.A(_10190_),
    .B(_10191_),
    .X(_02660_));
 sky130_fd_sc_hd__and2_1 _26859_ (.A(_10084_),
    .B(_10070_),
    .X(_10192_));
 sky130_fd_sc_hd__o21bai_4 _26860_ (.A1(_10068_),
    .A2(_10085_),
    .B1_N(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__a2bb2oi_4 _26861_ (.A1_N(_14368_),
    .A2_N(_10063_),
    .B1(_10062_),
    .B2(_10064_),
    .Y(_10194_));
 sky130_fd_sc_hd__a2bb2oi_4 _26862_ (.A1_N(_14385_),
    .A2_N(_10072_),
    .B1(_10071_),
    .B2(_10073_),
    .Y(_10195_));
 sky130_fd_sc_hd__and2_2 _26863_ (.A(_07106_),
    .B(_06279_),
    .X(_10196_));
 sky130_fd_sc_hd__nand3_4 _26864_ (.A(_08627_),
    .B(_08628_),
    .C(_06019_),
    .Y(_10197_));
 sky130_fd_sc_hd__a22o_2 _26865_ (.A1(_07262_),
    .A2(_08720_),
    .B1(_08405_),
    .B2(_07650_),
    .X(_10198_));
 sky130_fd_sc_hd__o21ai_4 _26866_ (.A1(_06034_),
    .A2(_10197_),
    .B1(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__xor2_4 _26867_ (.A(_10196_),
    .B(_10199_),
    .X(_10200_));
 sky130_fd_sc_hd__xnor2_4 _26868_ (.A(_10195_),
    .B(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__xnor2_4 _26869_ (.A(_10194_),
    .B(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__or2b_2 _26870_ (.A(_10082_),
    .B_N(_10077_),
    .X(_10203_));
 sky130_fd_sc_hd__o21ai_4 _26871_ (.A1(_10075_),
    .A2(_10083_),
    .B1(_10203_),
    .Y(_10204_));
 sky130_fd_sc_hd__and2_2 _26872_ (.A(_07873_),
    .B(_05770_),
    .X(_10205_));
 sky130_fd_sc_hd__nand3_4 _26873_ (.A(_08396_),
    .B(_09162_),
    .C(_06161_),
    .Y(_10206_));
 sky130_fd_sc_hd__a22o_2 _26874_ (.A1(_08636_),
    .A2(_05513_),
    .B1(_09162_),
    .B2(_05691_),
    .X(_10207_));
 sky130_fd_sc_hd__o21ai_4 _26875_ (.A1(_08210_),
    .A2(_10206_),
    .B1(_10207_),
    .Y(_10208_));
 sky130_fd_sc_hd__xor2_4 _26876_ (.A(_10205_),
    .B(_10208_),
    .X(_10209_));
 sky130_fd_sc_hd__nand3b_2 _26877_ (.A_N(_10079_),
    .B(_09876_),
    .C(_14405_),
    .Y(_10210_));
 sky130_fd_sc_hd__o31ai_4 _26878_ (.A1(_13967_),
    .A2(_05418_),
    .A3(_10081_),
    .B1(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__and2_2 _26879_ (.A(_09172_),
    .B(_08264_),
    .X(_10212_));
 sky130_fd_sc_hd__nand2_2 _26880_ (.A(_09174_),
    .B(_05321_),
    .Y(_10213_));
 sky130_fd_sc_hd__and2b_1 _26881_ (.A_N(_05613_),
    .B(_09176_),
    .X(_10214_));
 sky130_fd_sc_hd__xor2_4 _26882_ (.A(_10213_),
    .B(_10214_),
    .X(_10215_));
 sky130_fd_sc_hd__xor2_4 _26883_ (.A(_10212_),
    .B(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__xor2_4 _26884_ (.A(_10211_),
    .B(_10216_),
    .X(_10217_));
 sky130_fd_sc_hd__xor2_4 _26885_ (.A(_10209_),
    .B(_10217_),
    .X(_10218_));
 sky130_fd_sc_hd__xnor2_4 _26886_ (.A(_10204_),
    .B(_10218_),
    .Y(_10219_));
 sky130_fd_sc_hd__xor2_4 _26887_ (.A(_10202_),
    .B(_10219_),
    .X(_10220_));
 sky130_fd_sc_hd__nor2_4 _26888_ (.A(_10193_),
    .B(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__and2_1 _26889_ (.A(_10220_),
    .B(_10193_),
    .X(_10222_));
 sky130_fd_sc_hd__nor2_1 _26890_ (.A(_10051_),
    .B(_10052_),
    .Y(_10223_));
 sky130_fd_sc_hd__o21ba_2 _26891_ (.A1(_10046_),
    .A2(_10053_),
    .B1_N(_10223_),
    .X(_10224_));
 sky130_fd_sc_hd__nor2_1 _26892_ (.A(_10061_),
    .B(_10066_),
    .Y(_10225_));
 sky130_fd_sc_hd__o21bai_4 _26893_ (.A1(_10060_),
    .A2(_10067_),
    .B1_N(_10225_),
    .Y(_10226_));
 sky130_fd_sc_hd__and2_2 _26894_ (.A(_06059_),
    .B(_06957_),
    .X(_10227_));
 sky130_fd_sc_hd__nand3_4 _26895_ (.A(_08425_),
    .B(_09379_),
    .C(_08701_),
    .Y(_10228_));
 sky130_fd_sc_hd__a22o_2 _26896_ (.A1(_14010_),
    .A2(_07033_),
    .B1(_14015_),
    .B2(_07205_),
    .X(_10229_));
 sky130_fd_sc_hd__o21ai_4 _26897_ (.A1(_08699_),
    .A2(_10228_),
    .B1(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__xor2_4 _26898_ (.A(_10227_),
    .B(_10230_),
    .X(_10231_));
 sky130_fd_sc_hd__a2bb2oi_4 _26899_ (.A1_N(_14347_),
    .A2_N(_10048_),
    .B1(_10047_),
    .B2(_10049_),
    .Y(_10232_));
 sky130_fd_sc_hd__and2_2 _26900_ (.A(_06649_),
    .B(_06587_),
    .X(_10233_));
 sky130_fd_sc_hd__nand3_4 _26901_ (.A(_08431_),
    .B(_08432_),
    .C(_06165_),
    .Y(_10234_));
 sky130_fd_sc_hd__a22o_2 _26902_ (.A1(_08269_),
    .A2(_07648_),
    .B1(_06647_),
    .B2(_07046_),
    .X(_10235_));
 sky130_fd_sc_hd__o21ai_4 _26903_ (.A1(_14339_),
    .A2(_10234_),
    .B1(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__xor2_4 _26904_ (.A(_10233_),
    .B(_10236_),
    .X(_10237_));
 sky130_fd_sc_hd__xnor2_4 _26905_ (.A(_10232_),
    .B(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__xor2_4 _26906_ (.A(_10231_),
    .B(_10238_),
    .X(_10239_));
 sky130_fd_sc_hd__xnor2_4 _26907_ (.A(_10226_),
    .B(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__xor2_2 _26908_ (.A(_10224_),
    .B(_10240_),
    .X(_10241_));
 sky130_vsdinv _26909_ (.A(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__o21a_1 _26910_ (.A1(_10221_),
    .A2(_10222_),
    .B1(_10242_),
    .X(_10243_));
 sky130_fd_sc_hd__nand2_1 _26911_ (.A(_10220_),
    .B(_10193_),
    .Y(_10244_));
 sky130_fd_sc_hd__nor3b_4 _26912_ (.A(_10242_),
    .B(_10221_),
    .C_N(_10244_),
    .Y(_10245_));
 sky130_fd_sc_hd__and2_1 _26913_ (.A(_10086_),
    .B(_10059_),
    .X(_10246_));
 sky130_fd_sc_hd__o21bai_2 _26914_ (.A1(_10057_),
    .A2(_10087_),
    .B1_N(_10246_),
    .Y(_10247_));
 sky130_fd_sc_hd__o21bai_2 _26915_ (.A1(_10243_),
    .A2(_10245_),
    .B1_N(_10247_),
    .Y(_10248_));
 sky130_vsdinv _26916_ (.A(_10245_),
    .Y(_10249_));
 sky130_fd_sc_hd__nand3b_4 _26917_ (.A_N(_10243_),
    .B(_10247_),
    .C(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__or2b_1 _26918_ (.A(_10121_),
    .B_N(_10109_),
    .X(_10251_));
 sky130_fd_sc_hd__nand2_1 _26919_ (.A(_10120_),
    .B(_10111_),
    .Y(_10252_));
 sky130_fd_sc_hd__and2_1 _26920_ (.A(_10251_),
    .B(_10252_),
    .X(_10253_));
 sky130_fd_sc_hd__nand2_4 _26921_ (.A(_05445_),
    .B(\pcpi_mul.rs1[31] ),
    .Y(_10254_));
 sky130_fd_sc_hd__nand2_8 _26922_ (.A(_12776_),
    .B(_05271_),
    .Y(_10255_));
 sky130_fd_sc_hd__xnor2_4 _26923_ (.A(_10254_),
    .B(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__xor2_4 _26924_ (.A(_10104_),
    .B(_10256_),
    .X(_10257_));
 sky130_fd_sc_hd__a2bb2oi_4 _26925_ (.A1_N(_14292_),
    .A2_N(_10098_),
    .B1(_10097_),
    .B2(_10099_),
    .Y(_10258_));
 sky130_fd_sc_hd__and2_2 _26926_ (.A(_05441_),
    .B(_08078_),
    .X(_10259_));
 sky130_fd_sc_hd__nand3_4 _26927_ (.A(_07655_),
    .B(_14042_),
    .C(_07584_),
    .Y(_10260_));
 sky130_fd_sc_hd__a22o_2 _26928_ (.A1(_05955_),
    .A2(\pcpi_mul.rs1[28] ),
    .B1(_08199_),
    .B2(\pcpi_mul.rs1[29] ),
    .X(_10261_));
 sky130_fd_sc_hd__o21ai_4 _26929_ (.A1(_14285_),
    .A2(_10260_),
    .B1(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__xor2_4 _26930_ (.A(_10259_),
    .B(_10262_),
    .X(_10263_));
 sky130_fd_sc_hd__xnor2_4 _26931_ (.A(_10258_),
    .B(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__xor2_4 _26932_ (.A(_10257_),
    .B(_10264_),
    .X(_10265_));
 sky130_fd_sc_hd__nor2_1 _26933_ (.A(_10113_),
    .B(_10118_),
    .Y(_10266_));
 sky130_fd_sc_hd__o21bai_2 _26934_ (.A1(_10112_),
    .A2(_10119_),
    .B1_N(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__a2bb2oi_4 _26935_ (.A1_N(_14310_),
    .A2_N(_10115_),
    .B1(_10114_),
    .B2(_10116_),
    .Y(_10268_));
 sky130_fd_sc_hd__a2bb2oi_4 _26936_ (.A1_N(_14327_),
    .A2_N(_10043_),
    .B1(_10042_),
    .B2(_10044_),
    .Y(_10269_));
 sky130_fd_sc_hd__and2_2 _26937_ (.A(_06489_),
    .B(_08782_),
    .X(_10270_));
 sky130_fd_sc_hd__nand3_4 _26938_ (.A(_06349_),
    .B(_08357_),
    .C(_07209_),
    .Y(_10271_));
 sky130_fd_sc_hd__a22o_2 _26939_ (.A1(_06349_),
    .A2(_07786_),
    .B1(_14027_),
    .B2(\pcpi_mul.rs1[26] ),
    .X(_10272_));
 sky130_fd_sc_hd__o21ai_4 _26940_ (.A1(_14303_),
    .A2(_10271_),
    .B1(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__xor2_4 _26941_ (.A(_10270_),
    .B(_10273_),
    .X(_10274_));
 sky130_fd_sc_hd__xnor2_4 _26942_ (.A(_10269_),
    .B(_10274_),
    .Y(_10275_));
 sky130_fd_sc_hd__xor2_4 _26943_ (.A(_10268_),
    .B(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__xnor2_2 _26944_ (.A(_10267_),
    .B(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__xnor2_2 _26945_ (.A(_10265_),
    .B(_10277_),
    .Y(_10278_));
 sky130_fd_sc_hd__and2_1 _26946_ (.A(_10054_),
    .B(_10041_),
    .X(_10279_));
 sky130_fd_sc_hd__o21bai_4 _26947_ (.A1(_10039_),
    .A2(_10055_),
    .B1_N(_10279_),
    .Y(_10280_));
 sky130_fd_sc_hd__xor2_2 _26948_ (.A(_10278_),
    .B(_10280_),
    .X(_10281_));
 sky130_fd_sc_hd__xor2_1 _26949_ (.A(_10253_),
    .B(_10281_),
    .X(_10282_));
 sky130_fd_sc_hd__a21boi_1 _26950_ (.A1(_10248_),
    .A2(_10250_),
    .B1_N(_10282_),
    .Y(_10283_));
 sky130_vsdinv _26951_ (.A(_10283_),
    .Y(_10284_));
 sky130_fd_sc_hd__nand3b_4 _26952_ (.A_N(_10282_),
    .B(_10248_),
    .C(_10250_),
    .Y(_10285_));
 sky130_fd_sc_hd__nand2_2 _26953_ (.A(_10128_),
    .B(_10093_),
    .Y(_10286_));
 sky130_fd_sc_hd__a21o_1 _26954_ (.A1(_10284_),
    .A2(_10285_),
    .B1(_10286_),
    .X(_10287_));
 sky130_fd_sc_hd__nand3_4 _26955_ (.A(_10284_),
    .B(_10286_),
    .C(_10285_),
    .Y(_10288_));
 sky130_fd_sc_hd__nor2_2 _26956_ (.A(_10137_),
    .B(_10146_),
    .Y(_10289_));
 sky130_fd_sc_hd__a21oi_4 _26957_ (.A1(_10139_),
    .A2(_10145_),
    .B1(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__nand2_1 _26958_ (.A(_10143_),
    .B(_10135_),
    .Y(_10291_));
 sky130_fd_sc_hd__o21a_2 _26959_ (.A1(_10142_),
    .A2(_10144_),
    .B1(_10291_),
    .X(_10292_));
 sky130_fd_sc_hd__nor2_1 _26960_ (.A(_10096_),
    .B(_10101_),
    .Y(_10293_));
 sky130_fd_sc_hd__o21bai_4 _26961_ (.A1(_10102_),
    .A2(_10108_),
    .B1_N(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__inv_4 _26962_ (.A(_10104_),
    .Y(_10295_));
 sky130_fd_sc_hd__o21ai_4 _26963_ (.A1(_10295_),
    .A2(_10107_),
    .B1(_10105_),
    .Y(_10296_));
 sky130_fd_sc_hd__xnor2_4 _26964_ (.A(_09968_),
    .B(_10296_),
    .Y(_10297_));
 sky130_fd_sc_hd__xor2_4 _26965_ (.A(_10142_),
    .B(_10297_),
    .X(_10298_));
 sky130_fd_sc_hd__xnor2_4 _26966_ (.A(_10294_),
    .B(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__xor2_4 _26967_ (.A(_10292_),
    .B(_10299_),
    .X(_10300_));
 sky130_fd_sc_hd__xor2_4 _26968_ (.A(_10290_),
    .B(_10300_),
    .X(_10301_));
 sky130_fd_sc_hd__nor2_2 _26969_ (.A(_09985_),
    .B(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__and2_1 _26970_ (.A(_10301_),
    .B(_10149_),
    .X(_10303_));
 sky130_fd_sc_hd__or2b_1 _26971_ (.A(_10124_),
    .B_N(_10122_),
    .X(_10304_));
 sky130_fd_sc_hd__o21ai_2 _26972_ (.A1(_10095_),
    .A2(_10125_),
    .B1(_10304_),
    .Y(_10305_));
 sky130_fd_sc_hd__o21bai_2 _26973_ (.A1(_10302_),
    .A2(_10303_),
    .B1_N(_10305_),
    .Y(_10306_));
 sky130_vsdinv _26974_ (.A(_10302_),
    .Y(_10307_));
 sky130_fd_sc_hd__nand3b_4 _26975_ (.A_N(_10303_),
    .B(_10305_),
    .C(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__or2b_1 _26976_ (.A(_10134_),
    .B_N(_10147_),
    .X(_10309_));
 sky130_fd_sc_hd__o21a_1 _26977_ (.A1(_09985_),
    .A2(_10148_),
    .B1(_10309_),
    .X(_10310_));
 sky130_vsdinv _26978_ (.A(_10310_),
    .Y(_10311_));
 sky130_fd_sc_hd__a21o_1 _26979_ (.A1(_10306_),
    .A2(_10308_),
    .B1(_10311_),
    .X(_10312_));
 sky130_fd_sc_hd__nand3_4 _26980_ (.A(_10306_),
    .B(_10308_),
    .C(_10311_),
    .Y(_10313_));
 sky130_fd_sc_hd__nand2_4 _26981_ (.A(_10312_),
    .B(_10313_),
    .Y(_10314_));
 sky130_fd_sc_hd__a21boi_2 _26982_ (.A1(_10287_),
    .A2(_10288_),
    .B1_N(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__a21oi_4 _26983_ (.A1(_10284_),
    .A2(_10285_),
    .B1(_10286_),
    .Y(_10316_));
 sky130_fd_sc_hd__nor3b_4 _26984_ (.A(_10314_),
    .B(_10316_),
    .C_N(_10288_),
    .Y(_10317_));
 sky130_vsdinv _26985_ (.A(_10127_),
    .Y(_10318_));
 sky130_fd_sc_hd__a21oi_1 _26986_ (.A1(_10318_),
    .A2(_10128_),
    .B1(_10130_),
    .Y(_10319_));
 sky130_fd_sc_hd__o21ai_2 _26987_ (.A1(_10161_),
    .A2(_10319_),
    .B1(_10132_),
    .Y(_10320_));
 sky130_fd_sc_hd__o21bai_4 _26988_ (.A1(_10315_),
    .A2(_10317_),
    .B1_N(_10320_),
    .Y(_10321_));
 sky130_fd_sc_hd__a21bo_1 _26989_ (.A1(_10287_),
    .A2(_10288_),
    .B1_N(_10314_),
    .X(_10322_));
 sky130_fd_sc_hd__nand3b_2 _26990_ (.A_N(_10314_),
    .B(_10287_),
    .C(_10288_),
    .Y(_10323_));
 sky130_fd_sc_hd__nand3_4 _26991_ (.A(_10322_),
    .B(_10320_),
    .C(_10323_),
    .Y(_10324_));
 sky130_fd_sc_hd__buf_8 _26992_ (.A(_10000_),
    .X(_10325_));
 sky130_fd_sc_hd__a21oi_4 _26993_ (.A1(_10160_),
    .A2(_10156_),
    .B1(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__and3_1 _26994_ (.A(_10160_),
    .B(_10000_),
    .C(_10156_),
    .X(_10327_));
 sky130_fd_sc_hd__nor2_2 _26995_ (.A(_10326_),
    .B(_10327_),
    .Y(_10328_));
 sky130_fd_sc_hd__a21oi_1 _26996_ (.A1(_10321_),
    .A2(_10324_),
    .B1(_10328_),
    .Y(_10329_));
 sky130_fd_sc_hd__nand3_4 _26997_ (.A(_10321_),
    .B(_10328_),
    .C(_10324_),
    .Y(_10330_));
 sky130_vsdinv _26998_ (.A(_10330_),
    .Y(_10331_));
 sky130_vsdinv _26999_ (.A(_10172_),
    .Y(_10332_));
 sky130_fd_sc_hd__o21ai_2 _27000_ (.A1(_10332_),
    .A2(_10167_),
    .B1(_10168_),
    .Y(_10333_));
 sky130_fd_sc_hd__o21bai_2 _27001_ (.A1(_10329_),
    .A2(_10331_),
    .B1_N(_10333_),
    .Y(_10334_));
 sky130_fd_sc_hd__o2bb2ai_2 _27002_ (.A1_N(_10324_),
    .A2_N(_10321_),
    .B1(_10326_),
    .B2(_10327_),
    .Y(_10335_));
 sky130_fd_sc_hd__nand3_4 _27003_ (.A(_10335_),
    .B(_10333_),
    .C(_10330_),
    .Y(_10336_));
 sky130_fd_sc_hd__buf_4 _27004_ (.A(_10325_),
    .X(_10337_));
 sky130_fd_sc_hd__buf_8 _27005_ (.A(net413),
    .X(_10338_));
 sky130_fd_sc_hd__a21oi_4 _27006_ (.A1(_09989_),
    .A2(_09983_),
    .B1(_10338_),
    .Y(_10339_));
 sky130_fd_sc_hd__a21oi_1 _27007_ (.A1(_10334_),
    .A2(_10336_),
    .B1(_10339_),
    .Y(_10340_));
 sky130_fd_sc_hd__nand3_4 _27008_ (.A(_10334_),
    .B(_10339_),
    .C(_10336_),
    .Y(_10341_));
 sky130_vsdinv _27009_ (.A(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__o21ai_2 _27010_ (.A1(_10181_),
    .A2(_10182_),
    .B1(_10177_),
    .Y(_10343_));
 sky130_fd_sc_hd__o21bai_1 _27011_ (.A1(_10340_),
    .A2(_10342_),
    .B1_N(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__nand3b_4 _27012_ (.A_N(_10340_),
    .B(_10341_),
    .C(_10343_),
    .Y(_10345_));
 sky130_fd_sc_hd__nand2_2 _27013_ (.A(_10344_),
    .B(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__a21oi_1 _27014_ (.A1(_10187_),
    .A2(_10188_),
    .B1(_10185_),
    .Y(_10347_));
 sky130_fd_sc_hd__a21oi_2 _27015_ (.A1(_10025_),
    .A2(_10189_),
    .B1(_10347_),
    .Y(_10348_));
 sky130_fd_sc_hd__nor3_4 _27016_ (.A(_10026_),
    .B(_10190_),
    .C(_10037_),
    .Y(_10349_));
 sky130_fd_sc_hd__nor2_2 _27017_ (.A(_10348_),
    .B(_10349_),
    .Y(_10350_));
 sky130_fd_sc_hd__xor2_1 _27018_ (.A(_10346_),
    .B(_10350_),
    .X(_02661_));
 sky130_fd_sc_hd__nor2_1 _27019_ (.A(_10232_),
    .B(_10237_),
    .Y(_10351_));
 sky130_fd_sc_hd__o21ba_2 _27020_ (.A1(_10231_),
    .A2(_10238_),
    .B1_N(_10351_),
    .X(_10352_));
 sky130_fd_sc_hd__nor2_1 _27021_ (.A(_10195_),
    .B(_10200_),
    .Y(_10353_));
 sky130_fd_sc_hd__o21bai_4 _27022_ (.A1(_10194_),
    .A2(_10201_),
    .B1_N(_10353_),
    .Y(_10354_));
 sky130_fd_sc_hd__and2_2 _27023_ (.A(_08261_),
    .B(_07210_),
    .X(_10355_));
 sky130_fd_sc_hd__nand3_4 _27024_ (.A(_08660_),
    .B(_08426_),
    .C(_07206_),
    .Y(_10356_));
 sky130_fd_sc_hd__a22o_2 _27025_ (.A1(_06895_),
    .A2(_07036_),
    .B1(_06896_),
    .B2(_07039_),
    .X(_10357_));
 sky130_fd_sc_hd__o21ai_4 _27026_ (.A1(_14315_),
    .A2(_10356_),
    .B1(_10357_),
    .Y(_10358_));
 sky130_fd_sc_hd__xor2_4 _27027_ (.A(_10355_),
    .B(_10358_),
    .X(_10359_));
 sky130_fd_sc_hd__a2bb2oi_4 _27028_ (.A1_N(_14341_),
    .A2_N(_10234_),
    .B1(_10233_),
    .B2(_10235_),
    .Y(_10360_));
 sky130_fd_sc_hd__and2_2 _27029_ (.A(_06649_),
    .B(_06940_),
    .X(_10361_));
 sky130_fd_sc_hd__nand3_4 _27030_ (.A(_08667_),
    .B(_08864_),
    .C(_07746_),
    .Y(_10362_));
 sky130_fd_sc_hd__a22o_2 _27031_ (.A1(_07246_),
    .A2(_07046_),
    .B1(_08432_),
    .B2(_06760_),
    .X(_10363_));
 sky130_fd_sc_hd__o21ai_4 _27032_ (.A1(_14333_),
    .A2(_10362_),
    .B1(_10363_),
    .Y(_10364_));
 sky130_fd_sc_hd__xor2_4 _27033_ (.A(_10361_),
    .B(_10364_),
    .X(_10365_));
 sky130_fd_sc_hd__xnor2_4 _27034_ (.A(_10360_),
    .B(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__xor2_4 _27035_ (.A(_10359_),
    .B(_10366_),
    .X(_10367_));
 sky130_fd_sc_hd__xnor2_4 _27036_ (.A(_10354_),
    .B(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__xor2_2 _27037_ (.A(_10352_),
    .B(_10368_),
    .X(_10369_));
 sky130_vsdinv _27038_ (.A(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__and2_1 _27039_ (.A(_10218_),
    .B(_10204_),
    .X(_10371_));
 sky130_fd_sc_hd__o21bai_4 _27040_ (.A1(_10202_),
    .A2(_10219_),
    .B1_N(_10371_),
    .Y(_10372_));
 sky130_fd_sc_hd__a2bb2oi_4 _27041_ (.A1_N(_14361_),
    .A2_N(_10197_),
    .B1(_10196_),
    .B2(_10198_),
    .Y(_10373_));
 sky130_fd_sc_hd__a2bb2oi_4 _27042_ (.A1_N(_14379_),
    .A2_N(_10206_),
    .B1(_10205_),
    .B2(_10207_),
    .Y(_10374_));
 sky130_fd_sc_hd__nand2_2 _27043_ (.A(_08400_),
    .B(_06584_),
    .Y(_10375_));
 sky130_fd_sc_hd__or4_4 _27044_ (.A(_08402_),
    .B(_13989_),
    .C(_14352_),
    .D(_14359_),
    .X(_10376_));
 sky130_fd_sc_hd__a22o_1 _27045_ (.A1(_08404_),
    .A2(_07650_),
    .B1(_08405_),
    .B2(_06155_),
    .X(_10377_));
 sky130_fd_sc_hd__nand2_2 _27046_ (.A(_10376_),
    .B(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__xnor2_4 _27047_ (.A(_10375_),
    .B(_10378_),
    .Y(_10379_));
 sky130_fd_sc_hd__xnor2_4 _27048_ (.A(_10374_),
    .B(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__xnor2_4 _27049_ (.A(_10373_),
    .B(_10380_),
    .Y(_10381_));
 sky130_fd_sc_hd__or2b_1 _27050_ (.A(_10216_),
    .B_N(_10211_),
    .X(_10382_));
 sky130_fd_sc_hd__o21ai_4 _27051_ (.A1(_10209_),
    .A2(_10217_),
    .B1(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__and2_2 _27052_ (.A(_08634_),
    .B(_05778_),
    .X(_10384_));
 sky130_fd_sc_hd__nand3_4 _27053_ (.A(_08636_),
    .B(_08637_),
    .C(_05691_),
    .Y(_10385_));
 sky130_fd_sc_hd__a22o_2 _27054_ (.A1(_08374_),
    .A2(_09198_),
    .B1(_09164_),
    .B2(_05905_),
    .X(_10386_));
 sky130_fd_sc_hd__o21ai_4 _27055_ (.A1(_14372_),
    .A2(_10385_),
    .B1(_10386_),
    .Y(_10387_));
 sky130_fd_sc_hd__xor2_4 _27056_ (.A(_10384_),
    .B(_10387_),
    .X(_10388_));
 sky130_fd_sc_hd__nand3b_2 _27057_ (.A_N(_10213_),
    .B(_08526_),
    .C(_05874_),
    .Y(_10389_));
 sky130_fd_sc_hd__o31ai_4 _27058_ (.A1(_09168_),
    .A2(_07668_),
    .A3(_10215_),
    .B1(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__and2_2 _27059_ (.A(_08644_),
    .B(_05512_),
    .X(_10391_));
 sky130_fd_sc_hd__nand2_2 _27060_ (.A(_08646_),
    .B(_06002_),
    .Y(_10392_));
 sky130_fd_sc_hd__and2b_1 _27061_ (.A_N(_05882_),
    .B(_08383_),
    .X(_10393_));
 sky130_fd_sc_hd__xor2_4 _27062_ (.A(_10392_),
    .B(_10393_),
    .X(_10394_));
 sky130_fd_sc_hd__xor2_4 _27063_ (.A(_10391_),
    .B(_10394_),
    .X(_10395_));
 sky130_fd_sc_hd__xor2_4 _27064_ (.A(_10390_),
    .B(_10395_),
    .X(_10396_));
 sky130_fd_sc_hd__xor2_4 _27065_ (.A(_10388_),
    .B(_10396_),
    .X(_10397_));
 sky130_fd_sc_hd__xnor2_4 _27066_ (.A(_10383_),
    .B(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__xor2_4 _27067_ (.A(_10381_),
    .B(_10398_),
    .X(_10399_));
 sky130_fd_sc_hd__xnor2_1 _27068_ (.A(_10372_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__nor2_2 _27069_ (.A(_10370_),
    .B(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__and2_1 _27070_ (.A(_10400_),
    .B(_10370_),
    .X(_10402_));
 sky130_fd_sc_hd__o21ai_1 _27071_ (.A1(_10242_),
    .A2(_10221_),
    .B1(_10244_),
    .Y(_10403_));
 sky130_fd_sc_hd__o21ba_1 _27072_ (.A1(_10401_),
    .A2(_10402_),
    .B1_N(_10403_),
    .X(_10404_));
 sky130_vsdinv _27073_ (.A(_10404_),
    .Y(_10405_));
 sky130_fd_sc_hd__a211o_4 _27074_ (.A1(_10249_),
    .A2(_10244_),
    .B1(_10401_),
    .C1(_10402_),
    .X(_10406_));
 sky130_fd_sc_hd__or2b_1 _27075_ (.A(_10277_),
    .B_N(_10265_),
    .X(_10407_));
 sky130_fd_sc_hd__nand2_1 _27076_ (.A(_10276_),
    .B(_10267_),
    .Y(_10408_));
 sky130_fd_sc_hd__and2_2 _27077_ (.A(_10407_),
    .B(_10408_),
    .X(_10409_));
 sky130_fd_sc_hd__and2_1 _27078_ (.A(_10239_),
    .B(_10226_),
    .X(_10410_));
 sky130_fd_sc_hd__o21bai_4 _27079_ (.A1(_10224_),
    .A2(_10240_),
    .B1_N(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__nand2_4 _27080_ (.A(_12776_),
    .B(_14050_),
    .Y(_10412_));
 sky130_fd_sc_hd__xnor2_4 _27081_ (.A(_10255_),
    .B(_10412_),
    .Y(_10413_));
 sky130_fd_sc_hd__xor2_4 _27082_ (.A(_10295_),
    .B(_10413_),
    .X(_10414_));
 sky130_fd_sc_hd__clkinv_8 _27083_ (.A(_10414_),
    .Y(_10415_));
 sky130_fd_sc_hd__a2bb2oi_4 _27084_ (.A1_N(_08084_),
    .A2_N(_10260_),
    .B1(_10259_),
    .B2(_10261_),
    .Y(_10416_));
 sky130_fd_sc_hd__and2_2 _27085_ (.A(_05441_),
    .B(_08170_),
    .X(_10417_));
 sky130_fd_sc_hd__nand3_4 _27086_ (.A(_07281_),
    .B(_05531_),
    .C(_07784_),
    .Y(_10418_));
 sky130_fd_sc_hd__a22o_2 _27087_ (.A1(_14037_),
    .A2(_07784_),
    .B1(_14042_),
    .B2(_08077_),
    .X(_10419_));
 sky130_fd_sc_hd__o21ai_4 _27088_ (.A1(_14278_),
    .A2(_10418_),
    .B1(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__xor2_4 _27089_ (.A(_10417_),
    .B(_10420_),
    .X(_10421_));
 sky130_fd_sc_hd__xnor2_4 _27090_ (.A(_10416_),
    .B(_10421_),
    .Y(_10422_));
 sky130_fd_sc_hd__xor2_4 _27091_ (.A(_10415_),
    .B(_10422_),
    .X(_10423_));
 sky130_fd_sc_hd__nor2_1 _27092_ (.A(_10269_),
    .B(_10274_),
    .Y(_10424_));
 sky130_fd_sc_hd__o21bai_4 _27093_ (.A1(_10268_),
    .A2(_10275_),
    .B1_N(_10424_),
    .Y(_10425_));
 sky130_fd_sc_hd__a2bb2oi_4 _27094_ (.A1_N(_09222_),
    .A2_N(_10271_),
    .B1(_10270_),
    .B2(_10272_),
    .Y(_10426_));
 sky130_fd_sc_hd__a2bb2oi_4 _27095_ (.A1_N(_08699_),
    .A2_N(_10228_),
    .B1(_10227_),
    .B2(_10229_),
    .Y(_10427_));
 sky130_fd_sc_hd__and2_2 _27096_ (.A(_06355_),
    .B(_07584_),
    .X(_10428_));
 sky130_fd_sc_hd__nand3_4 _27097_ (.A(_08354_),
    .B(_08357_),
    .C(_07476_),
    .Y(_10429_));
 sky130_fd_sc_hd__a22o_2 _27098_ (.A1(_06349_),
    .A2(_07476_),
    .B1(_08357_),
    .B2(_07484_),
    .X(_10430_));
 sky130_fd_sc_hd__o21ai_4 _27099_ (.A1(_14296_),
    .A2(_10429_),
    .B1(_10430_),
    .Y(_10431_));
 sky130_fd_sc_hd__xor2_4 _27100_ (.A(_10428_),
    .B(_10431_),
    .X(_10432_));
 sky130_fd_sc_hd__xnor2_4 _27101_ (.A(_10427_),
    .B(_10432_),
    .Y(_10433_));
 sky130_fd_sc_hd__xor2_4 _27102_ (.A(_10426_),
    .B(_10433_),
    .X(_10434_));
 sky130_fd_sc_hd__xnor2_4 _27103_ (.A(_10425_),
    .B(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__xnor2_4 _27104_ (.A(_10423_),
    .B(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__xor2_4 _27105_ (.A(_10411_),
    .B(_10436_),
    .X(_10437_));
 sky130_fd_sc_hd__xor2_4 _27106_ (.A(_10409_),
    .B(_10437_),
    .X(_10438_));
 sky130_fd_sc_hd__a21boi_1 _27107_ (.A1(_10405_),
    .A2(_10406_),
    .B1_N(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__nand3b_4 _27108_ (.A_N(_10438_),
    .B(_10405_),
    .C(_10406_),
    .Y(_10440_));
 sky130_vsdinv _27109_ (.A(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__nand2_4 _27110_ (.A(_10285_),
    .B(_10250_),
    .Y(_10442_));
 sky130_fd_sc_hd__o21bai_2 _27111_ (.A1(_10439_),
    .A2(_10441_),
    .B1_N(_10442_),
    .Y(_10443_));
 sky130_fd_sc_hd__a21bo_2 _27112_ (.A1(_10405_),
    .A2(_10406_),
    .B1_N(_10438_),
    .X(_10444_));
 sky130_fd_sc_hd__nand3_4 _27113_ (.A(_10444_),
    .B(_10440_),
    .C(_10442_),
    .Y(_10445_));
 sky130_fd_sc_hd__clkbuf_4 _27114_ (.A(_10149_),
    .X(_10446_));
 sky130_fd_sc_hd__or2b_1 _27115_ (.A(_10290_),
    .B_N(_10300_),
    .X(_10447_));
 sky130_fd_sc_hd__o21a_2 _27116_ (.A1(_10446_),
    .A2(_10301_),
    .B1(_10447_),
    .X(_10448_));
 sky130_fd_sc_hd__nand2_1 _27117_ (.A(_10296_),
    .B(_10135_),
    .Y(_10449_));
 sky130_fd_sc_hd__o21a_2 _27118_ (.A1(_10142_),
    .A2(_10297_),
    .B1(_10449_),
    .X(_10450_));
 sky130_fd_sc_hd__nor2_1 _27119_ (.A(_10258_),
    .B(_10263_),
    .Y(_10451_));
 sky130_fd_sc_hd__o21bai_4 _27120_ (.A1(_10257_),
    .A2(_10264_),
    .B1_N(_10451_),
    .Y(_10452_));
 sky130_fd_sc_hd__nor2_1 _27121_ (.A(_10254_),
    .B(_10255_),
    .Y(_10453_));
 sky130_fd_sc_hd__o21bai_4 _27122_ (.A1(_10295_),
    .A2(_10256_),
    .B1_N(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__xnor2_4 _27123_ (.A(_10454_),
    .B(_09967_),
    .Y(_10455_));
 sky130_fd_sc_hd__xor2_4 _27124_ (.A(_10142_),
    .B(_10455_),
    .X(_10456_));
 sky130_fd_sc_hd__xnor2_4 _27125_ (.A(_10452_),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__xor2_4 _27126_ (.A(_10450_),
    .B(_10457_),
    .X(_10458_));
 sky130_fd_sc_hd__nor2_2 _27127_ (.A(_10292_),
    .B(_10299_),
    .Y(_10459_));
 sky130_fd_sc_hd__a21oi_4 _27128_ (.A1(_10294_),
    .A2(_10298_),
    .B1(_10459_),
    .Y(_10460_));
 sky130_fd_sc_hd__xor2_4 _27129_ (.A(_10458_),
    .B(_10460_),
    .X(_10461_));
 sky130_fd_sc_hd__and2_1 _27130_ (.A(_10461_),
    .B(_09793_),
    .X(_10462_));
 sky130_vsdinv _27131_ (.A(_10253_),
    .Y(_10463_));
 sky130_fd_sc_hd__and2_1 _27132_ (.A(_10280_),
    .B(_10278_),
    .X(_10464_));
 sky130_fd_sc_hd__a21o_1 _27133_ (.A1(_10281_),
    .A2(_10463_),
    .B1(_10464_),
    .X(_10465_));
 sky130_fd_sc_hd__nor2_1 _27134_ (.A(_10149_),
    .B(_10461_),
    .Y(_10466_));
 sky130_vsdinv _27135_ (.A(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__nand3b_4 _27136_ (.A_N(_10462_),
    .B(_10465_),
    .C(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__o21bai_2 _27137_ (.A1(_10466_),
    .A2(_10462_),
    .B1_N(_10465_),
    .Y(_10469_));
 sky130_fd_sc_hd__nand2_4 _27138_ (.A(_10468_),
    .B(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__xnor2_4 _27139_ (.A(_10448_),
    .B(_10470_),
    .Y(_10471_));
 sky130_vsdinv _27140_ (.A(_10471_),
    .Y(_10472_));
 sky130_fd_sc_hd__a21oi_1 _27141_ (.A1(_10443_),
    .A2(_10445_),
    .B1(_10472_),
    .Y(_10473_));
 sky130_fd_sc_hd__a21oi_4 _27142_ (.A1(_10444_),
    .A2(_10440_),
    .B1(_10442_),
    .Y(_10474_));
 sky130_vsdinv _27143_ (.A(_10445_),
    .Y(_10475_));
 sky130_fd_sc_hd__nor3_4 _27144_ (.A(_10471_),
    .B(_10474_),
    .C(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__o21ai_4 _27145_ (.A1(_10314_),
    .A2(_10316_),
    .B1(_10288_),
    .Y(_10477_));
 sky130_fd_sc_hd__o21bai_2 _27146_ (.A1(_10473_),
    .A2(_10476_),
    .B1_N(_10477_),
    .Y(_10478_));
 sky130_fd_sc_hd__nand2_1 _27147_ (.A(_10443_),
    .B(_10445_),
    .Y(_10479_));
 sky130_fd_sc_hd__nand2_2 _27148_ (.A(_10479_),
    .B(_10471_),
    .Y(_10480_));
 sky130_fd_sc_hd__nand3_4 _27149_ (.A(_10472_),
    .B(_10443_),
    .C(_10445_),
    .Y(_10481_));
 sky130_fd_sc_hd__nand3_4 _27150_ (.A(_10480_),
    .B(_10481_),
    .C(_10477_),
    .Y(_10482_));
 sky130_fd_sc_hd__nand2_1 _27151_ (.A(_10478_),
    .B(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__nand2_2 _27152_ (.A(_10313_),
    .B(_10308_),
    .Y(_10484_));
 sky130_fd_sc_hd__xor2_4 _27153_ (.A(net414),
    .B(_10484_),
    .X(_10485_));
 sky130_vsdinv _27154_ (.A(_10485_),
    .Y(_10486_));
 sky130_fd_sc_hd__nand2_2 _27155_ (.A(_10483_),
    .B(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__nand3_4 _27156_ (.A(_10478_),
    .B(_10485_),
    .C(_10482_),
    .Y(_10488_));
 sky130_fd_sc_hd__nand2_4 _27157_ (.A(_10330_),
    .B(_10324_),
    .Y(_10489_));
 sky130_fd_sc_hd__a21oi_4 _27158_ (.A1(_10487_),
    .A2(_10488_),
    .B1(_10489_),
    .Y(_10490_));
 sky130_fd_sc_hd__nand3_4 _27159_ (.A(_10487_),
    .B(_10488_),
    .C(_10489_),
    .Y(_10491_));
 sky130_vsdinv _27160_ (.A(_10491_),
    .Y(_10492_));
 sky130_fd_sc_hd__o21bai_2 _27161_ (.A1(_10490_),
    .A2(_10492_),
    .B1_N(_10326_),
    .Y(_10493_));
 sky130_fd_sc_hd__a21oi_1 _27162_ (.A1(_10478_),
    .A2(_10482_),
    .B1(_10485_),
    .Y(_10494_));
 sky130_fd_sc_hd__a21oi_4 _27163_ (.A1(_10480_),
    .A2(_10481_),
    .B1(_10477_),
    .Y(_10495_));
 sky130_vsdinv _27164_ (.A(_10482_),
    .Y(_10496_));
 sky130_fd_sc_hd__nor3_2 _27165_ (.A(_10486_),
    .B(_10495_),
    .C(_10496_),
    .Y(_10497_));
 sky130_fd_sc_hd__o21bai_1 _27166_ (.A1(_10494_),
    .A2(_10497_),
    .B1_N(_10489_),
    .Y(_10498_));
 sky130_fd_sc_hd__nand3_2 _27167_ (.A(_10498_),
    .B(_10326_),
    .C(_10491_),
    .Y(_10499_));
 sky130_fd_sc_hd__nand2_2 _27168_ (.A(_10341_),
    .B(_10336_),
    .Y(_10500_));
 sky130_fd_sc_hd__a21oi_2 _27169_ (.A1(_10493_),
    .A2(_10499_),
    .B1(_10500_),
    .Y(_10501_));
 sky130_fd_sc_hd__nand3_2 _27170_ (.A(_10493_),
    .B(_10500_),
    .C(_10499_),
    .Y(_10502_));
 sky130_vsdinv _27171_ (.A(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__nor2_2 _27172_ (.A(_10501_),
    .B(_10503_),
    .Y(_10504_));
 sky130_fd_sc_hd__o21ai_1 _27173_ (.A1(_10346_),
    .A2(_10350_),
    .B1(_10345_),
    .Y(_10505_));
 sky130_fd_sc_hd__xor2_1 _27174_ (.A(_10504_),
    .B(_10505_),
    .X(_02662_));
 sky130_fd_sc_hd__nor2_1 _27175_ (.A(_10360_),
    .B(_10365_),
    .Y(_10506_));
 sky130_fd_sc_hd__o21ba_2 _27176_ (.A1(_10359_),
    .A2(_10366_),
    .B1_N(_10506_),
    .X(_10507_));
 sky130_fd_sc_hd__and2_2 _27177_ (.A(_06060_),
    .B(_07569_),
    .X(_10508_));
 sky130_fd_sc_hd__nand3_4 _27178_ (.A(_08857_),
    .B(_08423_),
    .C(_07199_),
    .Y(_10509_));
 sky130_fd_sc_hd__a22o_2 _27179_ (.A1(_08660_),
    .A2(_08085_),
    .B1(_08859_),
    .B2(_07467_),
    .X(_10510_));
 sky130_fd_sc_hd__o21ai_4 _27180_ (.A1(_14310_),
    .A2(_10509_),
    .B1(_10510_),
    .Y(_10511_));
 sky130_fd_sc_hd__xor2_4 _27181_ (.A(_10508_),
    .B(_10511_),
    .X(_10512_));
 sky130_fd_sc_hd__a2bb2oi_4 _27182_ (.A1_N(_14335_),
    .A2_N(_10362_),
    .B1(_10361_),
    .B2(_10363_),
    .Y(_10513_));
 sky130_fd_sc_hd__and2_2 _27183_ (.A(_08673_),
    .B(_08330_),
    .X(_10514_));
 sky130_fd_sc_hd__buf_4 _27184_ (.A(_08667_),
    .X(_10515_));
 sky130_fd_sc_hd__clkbuf_4 _27185_ (.A(_08668_),
    .X(_10516_));
 sky130_fd_sc_hd__nand3_4 _27186_ (.A(_10515_),
    .B(_10516_),
    .C(_06761_),
    .Y(_10517_));
 sky130_fd_sc_hd__a22o_2 _27187_ (.A1(_07247_),
    .A2(_06761_),
    .B1(_09723_),
    .B2(_08701_),
    .X(_10518_));
 sky130_fd_sc_hd__o21ai_4 _27188_ (.A1(_14328_),
    .A2(_10517_),
    .B1(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__xor2_4 _27189_ (.A(_10514_),
    .B(_10519_),
    .X(_10520_));
 sky130_fd_sc_hd__xnor2_4 _27190_ (.A(_10513_),
    .B(_10520_),
    .Y(_10521_));
 sky130_fd_sc_hd__xor2_4 _27191_ (.A(_10512_),
    .B(_10521_),
    .X(_10522_));
 sky130_fd_sc_hd__nor2_1 _27192_ (.A(_10374_),
    .B(_10379_),
    .Y(_10523_));
 sky130_fd_sc_hd__o21bai_4 _27193_ (.A1(_10373_),
    .A2(_10380_),
    .B1_N(_10523_),
    .Y(_10524_));
 sky130_fd_sc_hd__xnor2_2 _27194_ (.A(_10522_),
    .B(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__xor2_1 _27195_ (.A(_10507_),
    .B(_10525_),
    .X(_10526_));
 sky130_fd_sc_hd__and2_1 _27196_ (.A(_10397_),
    .B(_10383_),
    .X(_10527_));
 sky130_fd_sc_hd__o21bai_2 _27197_ (.A1(_10381_),
    .A2(_10398_),
    .B1_N(_10527_),
    .Y(_10528_));
 sky130_fd_sc_hd__o21a_2 _27198_ (.A1(_10375_),
    .A2(_10378_),
    .B1(_10376_),
    .X(_10529_));
 sky130_fd_sc_hd__a2bb2oi_4 _27199_ (.A1_N(_14374_),
    .A2_N(_10385_),
    .B1(_10384_),
    .B2(_10386_),
    .Y(_10530_));
 sky130_fd_sc_hd__and2_2 _27200_ (.A(_08400_),
    .B(_07747_),
    .X(_10531_));
 sky130_fd_sc_hd__nand3_4 _27201_ (.A(_09152_),
    .B(_09153_),
    .C(_06279_),
    .Y(_10532_));
 sky130_fd_sc_hd__a22o_2 _27202_ (.A1(_08627_),
    .A2(_06155_),
    .B1(_08628_),
    .B2(_06431_),
    .X(_10533_));
 sky130_fd_sc_hd__o21ai_4 _27203_ (.A1(_14347_),
    .A2(_10532_),
    .B1(_10533_),
    .Y(_10534_));
 sky130_fd_sc_hd__xor2_4 _27204_ (.A(_10531_),
    .B(_10534_),
    .X(_10535_));
 sky130_fd_sc_hd__xnor2_4 _27205_ (.A(_10530_),
    .B(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__xnor2_4 _27206_ (.A(_10529_),
    .B(_10536_),
    .Y(_10537_));
 sky130_fd_sc_hd__or2b_1 _27207_ (.A(_10395_),
    .B_N(_10390_),
    .X(_10538_));
 sky130_fd_sc_hd__o21ai_4 _27208_ (.A1(_10388_),
    .A2(_10396_),
    .B1(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__and2_2 _27209_ (.A(_07873_),
    .B(_06147_),
    .X(_10540_));
 sky130_fd_sc_hd__nand3_4 _27210_ (.A(_09357_),
    .B(_08637_),
    .C(_05905_),
    .Y(_10541_));
 sky130_fd_sc_hd__a22o_2 _27211_ (.A1(_08636_),
    .A2(_05905_),
    .B1(_09164_),
    .B2(_06019_),
    .X(_10542_));
 sky130_fd_sc_hd__o21ai_4 _27212_ (.A1(_14366_),
    .A2(_10541_),
    .B1(_10542_),
    .Y(_10543_));
 sky130_fd_sc_hd__xor2_4 _27213_ (.A(_10540_),
    .B(_10543_),
    .X(_10544_));
 sky130_fd_sc_hd__nand3b_4 _27214_ (.A_N(_10392_),
    .B(_09169_),
    .C(_14394_),
    .Y(_10545_));
 sky130_fd_sc_hd__o31ai_4 _27215_ (.A1(_09168_),
    .A2(_14384_),
    .A3(_10394_),
    .B1(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__and2_2 _27216_ (.A(_09172_),
    .B(_09198_),
    .X(_10547_));
 sky130_fd_sc_hd__nand2_2 _27217_ (.A(_09174_),
    .B(_05915_),
    .Y(_10548_));
 sky130_fd_sc_hd__and2b_1 _27218_ (.A_N(_06002_),
    .B(_09176_),
    .X(_10549_));
 sky130_fd_sc_hd__xor2_4 _27219_ (.A(_10548_),
    .B(_10549_),
    .X(_10550_));
 sky130_fd_sc_hd__xor2_4 _27220_ (.A(_10547_),
    .B(_10550_),
    .X(_10551_));
 sky130_fd_sc_hd__xor2_4 _27221_ (.A(_10546_),
    .B(_10551_),
    .X(_10552_));
 sky130_fd_sc_hd__xor2_4 _27222_ (.A(_10544_),
    .B(_10552_),
    .X(_10553_));
 sky130_fd_sc_hd__xnor2_4 _27223_ (.A(_10539_),
    .B(_10553_),
    .Y(_10554_));
 sky130_fd_sc_hd__xor2_2 _27224_ (.A(_10537_),
    .B(_10554_),
    .X(_10555_));
 sky130_fd_sc_hd__xnor2_1 _27225_ (.A(_10528_),
    .B(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__or2b_2 _27226_ (.A(_10526_),
    .B_N(_10556_),
    .X(_10557_));
 sky130_fd_sc_hd__or2b_4 _27227_ (.A(_10556_),
    .B_N(_10526_),
    .X(_10558_));
 sky130_fd_sc_hd__a21o_1 _27228_ (.A1(_10399_),
    .A2(_10372_),
    .B1(_10401_),
    .X(_10559_));
 sky130_fd_sc_hd__a21o_2 _27229_ (.A1(_10557_),
    .A2(_10558_),
    .B1(_10559_),
    .X(_10560_));
 sky130_fd_sc_hd__nand3_4 _27230_ (.A(_10559_),
    .B(_10557_),
    .C(_10558_),
    .Y(_10561_));
 sky130_fd_sc_hd__or2b_1 _27231_ (.A(_10435_),
    .B_N(_10423_),
    .X(_10562_));
 sky130_fd_sc_hd__nand2_1 _27232_ (.A(_10434_),
    .B(_10425_),
    .Y(_10563_));
 sky130_fd_sc_hd__and2_1 _27233_ (.A(_10562_),
    .B(_10563_),
    .X(_10564_));
 sky130_fd_sc_hd__and2_1 _27234_ (.A(_10367_),
    .B(_10354_),
    .X(_10565_));
 sky130_fd_sc_hd__o21bai_4 _27235_ (.A1(_10352_),
    .A2(_10368_),
    .B1_N(_10565_),
    .Y(_10566_));
 sky130_fd_sc_hd__a2bb2oi_4 _27236_ (.A1_N(_14280_),
    .A2_N(_10418_),
    .B1(_10417_),
    .B2(_10419_),
    .Y(_10567_));
 sky130_fd_sc_hd__nand2_8 _27237_ (.A(_12778_),
    .B(_08710_),
    .Y(_10568_));
 sky130_fd_sc_hd__nand3_4 _27238_ (.A(_05956_),
    .B(_09071_),
    .C(_08078_),
    .Y(_10569_));
 sky130_fd_sc_hd__a22o_1 _27239_ (.A1(_07281_),
    .A2(_08077_),
    .B1(_05531_),
    .B2(_08170_),
    .X(_10570_));
 sky130_fd_sc_hd__o21ai_4 _27240_ (.A1(_14275_),
    .A2(_10569_),
    .B1(_10570_),
    .Y(_10571_));
 sky130_fd_sc_hd__xnor2_4 _27241_ (.A(_10568_),
    .B(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__xnor2_4 _27242_ (.A(_10567_),
    .B(_10572_),
    .Y(_10573_));
 sky130_fd_sc_hd__xor2_4 _27243_ (.A(_10415_),
    .B(_10573_),
    .X(_10574_));
 sky130_fd_sc_hd__nor2_1 _27244_ (.A(_10427_),
    .B(_10432_),
    .Y(_10575_));
 sky130_fd_sc_hd__o21bai_4 _27245_ (.A1(_10426_),
    .A2(_10433_),
    .B1_N(_10575_),
    .Y(_10576_));
 sky130_fd_sc_hd__a2bb2oi_4 _27246_ (.A1_N(_14299_),
    .A2_N(_10429_),
    .B1(_10428_),
    .B2(_10430_),
    .Y(_10577_));
 sky130_fd_sc_hd__a2bb2oi_4 _27247_ (.A1_N(_14315_),
    .A2_N(_10356_),
    .B1(_10355_),
    .B2(_10357_),
    .Y(_10578_));
 sky130_fd_sc_hd__and2_2 _27248_ (.A(_06355_),
    .B(_07784_),
    .X(_10579_));
 sky130_fd_sc_hd__nand3_4 _27249_ (.A(_06067_),
    .B(_06071_),
    .C(_08782_),
    .Y(_10580_));
 sky130_fd_sc_hd__a22o_2 _27250_ (.A1(_08354_),
    .A2(_07484_),
    .B1(_08355_),
    .B2(\pcpi_mul.rs1[28] ),
    .X(_10581_));
 sky130_fd_sc_hd__o21ai_4 _27251_ (.A1(_14290_),
    .A2(_10580_),
    .B1(_10581_),
    .Y(_10582_));
 sky130_fd_sc_hd__xor2_4 _27252_ (.A(_10579_),
    .B(_10582_),
    .X(_10583_));
 sky130_fd_sc_hd__xnor2_4 _27253_ (.A(_10578_),
    .B(_10583_),
    .Y(_10584_));
 sky130_fd_sc_hd__xor2_4 _27254_ (.A(_10577_),
    .B(_10584_),
    .X(_10585_));
 sky130_fd_sc_hd__xnor2_2 _27255_ (.A(_10576_),
    .B(_10585_),
    .Y(_10586_));
 sky130_fd_sc_hd__xnor2_2 _27256_ (.A(_10574_),
    .B(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__nor2_2 _27257_ (.A(_10566_),
    .B(_10587_),
    .Y(_10588_));
 sky130_fd_sc_hd__nand2_2 _27258_ (.A(_10587_),
    .B(_10566_),
    .Y(_10589_));
 sky130_fd_sc_hd__nor3b_4 _27259_ (.A(_10564_),
    .B(_10588_),
    .C_N(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__and2_1 _27260_ (.A(_10587_),
    .B(_10566_),
    .X(_10591_));
 sky130_fd_sc_hd__o21a_2 _27261_ (.A1(_10588_),
    .A2(_10591_),
    .B1(_10564_),
    .X(_10592_));
 sky130_fd_sc_hd__nor2_4 _27262_ (.A(_10590_),
    .B(_10592_),
    .Y(_10593_));
 sky130_fd_sc_hd__a21oi_2 _27263_ (.A1(_10560_),
    .A2(_10561_),
    .B1(_10593_),
    .Y(_10594_));
 sky130_fd_sc_hd__nand3_4 _27264_ (.A(_10560_),
    .B(_10593_),
    .C(_10561_),
    .Y(_10595_));
 sky130_vsdinv _27265_ (.A(_10595_),
    .Y(_10596_));
 sky130_fd_sc_hd__o21ai_4 _27266_ (.A1(_10438_),
    .A2(_10404_),
    .B1(_10406_),
    .Y(_10597_));
 sky130_fd_sc_hd__o21bai_4 _27267_ (.A1(_10594_),
    .A2(_10596_),
    .B1_N(_10597_),
    .Y(_10598_));
 sky130_fd_sc_hd__o2bb2ai_4 _27268_ (.A1_N(_10561_),
    .A2_N(_10560_),
    .B1(_10590_),
    .B2(_10592_),
    .Y(_10599_));
 sky130_fd_sc_hd__nand3_4 _27269_ (.A(_10599_),
    .B(_10595_),
    .C(_10597_),
    .Y(_10600_));
 sky130_fd_sc_hd__or2b_1 _27270_ (.A(_10460_),
    .B_N(_10458_),
    .X(_10601_));
 sky130_fd_sc_hd__o21a_4 _27271_ (.A1(_10446_),
    .A2(_10461_),
    .B1(_10601_),
    .X(_10602_));
 sky130_fd_sc_hd__nor2_2 _27272_ (.A(_10450_),
    .B(_10457_),
    .Y(_10603_));
 sky130_fd_sc_hd__a21oi_4 _27273_ (.A1(_10452_),
    .A2(_10456_),
    .B1(_10603_),
    .Y(_10604_));
 sky130_fd_sc_hd__nand2_1 _27274_ (.A(_10135_),
    .B(_10454_),
    .Y(_10605_));
 sky130_fd_sc_hd__o21a_2 _27275_ (.A1(_10142_),
    .A2(_10455_),
    .B1(_10605_),
    .X(_10606_));
 sky130_fd_sc_hd__nor2_1 _27276_ (.A(_10416_),
    .B(_10421_),
    .Y(_10607_));
 sky130_fd_sc_hd__o21bai_4 _27277_ (.A1(_10415_),
    .A2(_10422_),
    .B1_N(_10607_),
    .Y(_10608_));
 sky130_fd_sc_hd__inv_4 _27278_ (.A(_10141_),
    .Y(_10609_));
 sky130_fd_sc_hd__o22ai_4 _27279_ (.A1(_14051_),
    .A2(_10255_),
    .B1(_10295_),
    .B2(_10413_),
    .Y(_10610_));
 sky130_fd_sc_hd__xor2_4 _27280_ (.A(_10610_),
    .B(_09967_),
    .X(_10611_));
 sky130_fd_sc_hd__xor2_4 _27281_ (.A(_10609_),
    .B(_10611_),
    .X(_10612_));
 sky130_fd_sc_hd__xnor2_4 _27282_ (.A(_10608_),
    .B(_10612_),
    .Y(_10613_));
 sky130_fd_sc_hd__xor2_4 _27283_ (.A(_10606_),
    .B(_10613_),
    .X(_10614_));
 sky130_fd_sc_hd__xor2_2 _27284_ (.A(_10604_),
    .B(_10614_),
    .X(_10615_));
 sky130_fd_sc_hd__and2_1 _27285_ (.A(_10615_),
    .B(_09792_),
    .X(_10616_));
 sky130_vsdinv _27286_ (.A(_10409_),
    .Y(_10617_));
 sky130_fd_sc_hd__and2_1 _27287_ (.A(_10436_),
    .B(_10411_),
    .X(_10618_));
 sky130_fd_sc_hd__a21o_1 _27288_ (.A1(_10437_),
    .A2(_10617_),
    .B1(_10618_),
    .X(_10619_));
 sky130_fd_sc_hd__nor2_1 _27289_ (.A(_09793_),
    .B(_10615_),
    .Y(_10620_));
 sky130_vsdinv _27290_ (.A(_10620_),
    .Y(_10621_));
 sky130_fd_sc_hd__nand3b_4 _27291_ (.A_N(_10616_),
    .B(_10619_),
    .C(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__o21bai_2 _27292_ (.A1(_10620_),
    .A2(_10616_),
    .B1_N(_10619_),
    .Y(_10623_));
 sky130_fd_sc_hd__nand2_4 _27293_ (.A(_10622_),
    .B(_10623_),
    .Y(_10624_));
 sky130_fd_sc_hd__xor2_4 _27294_ (.A(_10602_),
    .B(_10624_),
    .X(_10625_));
 sky130_fd_sc_hd__a21o_1 _27295_ (.A1(_10598_),
    .A2(_10600_),
    .B1(_10625_),
    .X(_10626_));
 sky130_fd_sc_hd__nand3_4 _27296_ (.A(_10598_),
    .B(_10625_),
    .C(_10600_),
    .Y(_10627_));
 sky130_fd_sc_hd__o21ai_2 _27297_ (.A1(_10471_),
    .A2(_10474_),
    .B1(_10445_),
    .Y(_10628_));
 sky130_fd_sc_hd__nand3_4 _27298_ (.A(_10626_),
    .B(_10627_),
    .C(_10628_),
    .Y(_10629_));
 sky130_fd_sc_hd__a21oi_2 _27299_ (.A1(_10598_),
    .A2(_10600_),
    .B1(_10625_),
    .Y(_10630_));
 sky130_vsdinv _27300_ (.A(_10627_),
    .Y(_10631_));
 sky130_fd_sc_hd__o21bai_4 _27301_ (.A1(_10630_),
    .A2(_10631_),
    .B1_N(_10628_),
    .Y(_10632_));
 sky130_fd_sc_hd__o21a_2 _27302_ (.A1(_10448_),
    .A2(_10470_),
    .B1(_10468_),
    .X(_10633_));
 sky130_fd_sc_hd__nor2_8 _27303_ (.A(_10325_),
    .B(_10633_),
    .Y(_10634_));
 sky130_fd_sc_hd__o211a_2 _27304_ (.A1(_10448_),
    .A2(_10470_),
    .B1(_10000_),
    .C1(_10468_),
    .X(_10635_));
 sky130_fd_sc_hd__o2bb2ai_4 _27305_ (.A1_N(_10629_),
    .A2_N(_10632_),
    .B1(_10634_),
    .B2(_10635_),
    .Y(_10636_));
 sky130_fd_sc_hd__nor2_4 _27306_ (.A(_10635_),
    .B(_10634_),
    .Y(_10637_));
 sky130_fd_sc_hd__nand3_4 _27307_ (.A(_10632_),
    .B(_10637_),
    .C(_10629_),
    .Y(_10638_));
 sky130_fd_sc_hd__o21ai_4 _27308_ (.A1(_10486_),
    .A2(_10495_),
    .B1(_10482_),
    .Y(_10639_));
 sky130_fd_sc_hd__a21oi_4 _27309_ (.A1(_10636_),
    .A2(_10638_),
    .B1(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__nand3_4 _27310_ (.A(_10636_),
    .B(_10638_),
    .C(_10639_),
    .Y(_10641_));
 sky130_vsdinv _27311_ (.A(_10641_),
    .Y(_10642_));
 sky130_fd_sc_hd__a21oi_4 _27312_ (.A1(_10313_),
    .A2(_10308_),
    .B1(_10338_),
    .Y(_10643_));
 sky130_fd_sc_hd__o21bai_2 _27313_ (.A1(_10640_),
    .A2(_10642_),
    .B1_N(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__a21oi_1 _27314_ (.A1(_10632_),
    .A2(_10629_),
    .B1(_10637_),
    .Y(_10645_));
 sky130_vsdinv _27315_ (.A(_10638_),
    .Y(_10646_));
 sky130_fd_sc_hd__o21bai_2 _27316_ (.A1(_10645_),
    .A2(_10646_),
    .B1_N(_10639_),
    .Y(_10647_));
 sky130_fd_sc_hd__nand3_4 _27317_ (.A(_10647_),
    .B(_10643_),
    .C(_10641_),
    .Y(_10648_));
 sky130_vsdinv _27318_ (.A(_10326_),
    .Y(_10649_));
 sky130_fd_sc_hd__o21ai_4 _27319_ (.A1(_10649_),
    .A2(_10490_),
    .B1(_10491_),
    .Y(_10650_));
 sky130_fd_sc_hd__a21oi_2 _27320_ (.A1(_10644_),
    .A2(_10648_),
    .B1(_10650_),
    .Y(_10651_));
 sky130_fd_sc_hd__nand3_4 _27321_ (.A(_10644_),
    .B(_10648_),
    .C(_10650_),
    .Y(_10652_));
 sky130_vsdinv _27322_ (.A(_10652_),
    .Y(_10653_));
 sky130_fd_sc_hd__nor2_4 _27323_ (.A(_10651_),
    .B(_10653_),
    .Y(_10654_));
 sky130_fd_sc_hd__nor2_1 _27324_ (.A(_10026_),
    .B(_10190_),
    .Y(_10655_));
 sky130_fd_sc_hd__a21oi_1 _27325_ (.A1(_10498_),
    .A2(_10491_),
    .B1(_10326_),
    .Y(_10656_));
 sky130_fd_sc_hd__nor3_2 _27326_ (.A(_10649_),
    .B(_10490_),
    .C(_10492_),
    .Y(_10657_));
 sky130_fd_sc_hd__o21bai_1 _27327_ (.A1(_10656_),
    .A2(_10657_),
    .B1_N(_10500_),
    .Y(_10658_));
 sky130_fd_sc_hd__nand2_1 _27328_ (.A(_10658_),
    .B(_10502_),
    .Y(_10659_));
 sky130_fd_sc_hd__nor2_1 _27329_ (.A(_10346_),
    .B(_10659_),
    .Y(_10660_));
 sky130_fd_sc_hd__nand2_2 _27330_ (.A(_10655_),
    .B(_10660_),
    .Y(_10661_));
 sky130_vsdinv _27331_ (.A(_10346_),
    .Y(_10662_));
 sky130_fd_sc_hd__nand3_1 _27332_ (.A(_10504_),
    .B(_10662_),
    .C(_10348_),
    .Y(_10663_));
 sky130_fd_sc_hd__o21a_1 _27333_ (.A1(_10345_),
    .A2(_10501_),
    .B1(_10502_),
    .X(_10664_));
 sky130_fd_sc_hd__nand2_2 _27334_ (.A(_10663_),
    .B(_10664_),
    .Y(_10665_));
 sky130_fd_sc_hd__o21bai_4 _27335_ (.A1(_10661_),
    .A2(_10037_),
    .B1_N(_10665_),
    .Y(_10666_));
 sky130_fd_sc_hd__xor2_2 _27336_ (.A(_10654_),
    .B(_10666_),
    .X(_02663_));
 sky130_fd_sc_hd__and2_1 _27337_ (.A(_10553_),
    .B(_10539_),
    .X(_10667_));
 sky130_fd_sc_hd__o21bai_4 _27338_ (.A1(_10537_),
    .A2(_10554_),
    .B1_N(_10667_),
    .Y(_10668_));
 sky130_fd_sc_hd__a2bb2oi_4 _27339_ (.A1_N(_14348_),
    .A2_N(_10532_),
    .B1(_10531_),
    .B2(_10533_),
    .Y(_10669_));
 sky130_fd_sc_hd__a2bb2oi_4 _27340_ (.A1_N(_14368_),
    .A2_N(_10541_),
    .B1(_10540_),
    .B2(_10542_),
    .Y(_10670_));
 sky130_fd_sc_hd__and2_4 _27341_ (.A(_06888_),
    .B(_07481_),
    .X(_10671_));
 sky130_fd_sc_hd__buf_4 _27342_ (.A(_08404_),
    .X(_10672_));
 sky130_fd_sc_hd__nand3_4 _27343_ (.A(_10672_),
    .B(_07103_),
    .C(_08342_),
    .Y(_10673_));
 sky130_fd_sc_hd__a22o_2 _27344_ (.A1(_09152_),
    .A2(_06431_),
    .B1(_09153_),
    .B2(_06441_),
    .X(_10674_));
 sky130_fd_sc_hd__o21ai_4 _27345_ (.A1(_14340_),
    .A2(_10673_),
    .B1(_10674_),
    .Y(_10675_));
 sky130_fd_sc_hd__xor2_4 _27346_ (.A(_10671_),
    .B(_10675_),
    .X(_10676_));
 sky130_fd_sc_hd__xnor2_4 _27347_ (.A(_10670_),
    .B(_10676_),
    .Y(_10677_));
 sky130_fd_sc_hd__xnor2_4 _27348_ (.A(_10669_),
    .B(_10677_),
    .Y(_10678_));
 sky130_fd_sc_hd__or2b_1 _27349_ (.A(_10551_),
    .B_N(_10546_),
    .X(_10679_));
 sky130_fd_sc_hd__o21ai_4 _27350_ (.A1(_10544_),
    .A2(_10552_),
    .B1(_10679_),
    .Y(_10680_));
 sky130_fd_sc_hd__and2_2 _27351_ (.A(_07359_),
    .B(_06280_),
    .X(_10681_));
 sky130_fd_sc_hd__nand3_4 _27352_ (.A(_13972_),
    .B(_13978_),
    .C(_06020_),
    .Y(_10682_));
 sky130_fd_sc_hd__a22o_2 _27353_ (.A1(_08396_),
    .A2(_05778_),
    .B1(_13978_),
    .B2(_06285_),
    .X(_10683_));
 sky130_fd_sc_hd__o21ai_4 _27354_ (.A1(_14360_),
    .A2(_10682_),
    .B1(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__xor2_4 _27355_ (.A(_10681_),
    .B(_10684_),
    .X(_10685_));
 sky130_fd_sc_hd__nand3b_4 _27356_ (.A_N(_10548_),
    .B(_09876_),
    .C(_07668_),
    .Y(_10686_));
 sky130_fd_sc_hd__o31ai_4 _27357_ (.A1(_13967_),
    .A2(_08210_),
    .A3(_10550_),
    .B1(_10686_),
    .Y(_10687_));
 sky130_fd_sc_hd__and2_2 _27358_ (.A(_07945_),
    .B(_05769_),
    .X(_10688_));
 sky130_fd_sc_hd__nand2_2 _27359_ (.A(_13961_),
    .B(_05610_),
    .Y(_10689_));
 sky130_fd_sc_hd__and2b_1 _27360_ (.A_N(_05512_),
    .B(_12804_),
    .X(_10690_));
 sky130_fd_sc_hd__xor2_4 _27361_ (.A(_10689_),
    .B(_10690_),
    .X(_10691_));
 sky130_fd_sc_hd__xor2_4 _27362_ (.A(_10688_),
    .B(_10691_),
    .X(_10692_));
 sky130_fd_sc_hd__xor2_4 _27363_ (.A(_10687_),
    .B(_10692_),
    .X(_10693_));
 sky130_fd_sc_hd__xor2_4 _27364_ (.A(_10685_),
    .B(_10693_),
    .X(_10694_));
 sky130_fd_sc_hd__xnor2_4 _27365_ (.A(_10680_),
    .B(_10694_),
    .Y(_10695_));
 sky130_fd_sc_hd__xor2_4 _27366_ (.A(_10678_),
    .B(_10695_),
    .X(_10696_));
 sky130_fd_sc_hd__nor2_2 _27367_ (.A(_10668_),
    .B(_10696_),
    .Y(_10697_));
 sky130_fd_sc_hd__nand2_2 _27368_ (.A(_10696_),
    .B(_10668_),
    .Y(_10698_));
 sky130_vsdinv _27369_ (.A(_10698_),
    .Y(_10699_));
 sky130_fd_sc_hd__nor2_1 _27370_ (.A(_10513_),
    .B(_10520_),
    .Y(_10700_));
 sky130_fd_sc_hd__o21ba_4 _27371_ (.A1(_10512_),
    .A2(_10521_),
    .B1_N(_10700_),
    .X(_10701_));
 sky130_fd_sc_hd__nor2_1 _27372_ (.A(_10530_),
    .B(_10535_),
    .Y(_10702_));
 sky130_fd_sc_hd__o21bai_4 _27373_ (.A1(_10529_),
    .A2(_10536_),
    .B1_N(_10702_),
    .Y(_10703_));
 sky130_fd_sc_hd__and2_2 _27374_ (.A(_06060_),
    .B(_08070_),
    .X(_10704_));
 sky130_fd_sc_hd__clkbuf_4 _27375_ (.A(_09379_),
    .X(_10705_));
 sky130_fd_sc_hd__nand3_4 _27376_ (.A(_08857_),
    .B(_10705_),
    .C(_07468_),
    .Y(_10706_));
 sky130_fd_sc_hd__a22o_2 _27377_ (.A1(_08422_),
    .A2(_08885_),
    .B1(_08423_),
    .B2(_07775_),
    .X(_10707_));
 sky130_fd_sc_hd__o21ai_4 _27378_ (.A1(_09222_),
    .A2(_10706_),
    .B1(_10707_),
    .Y(_10708_));
 sky130_fd_sc_hd__xor2_4 _27379_ (.A(_10704_),
    .B(_10708_),
    .X(_10709_));
 sky130_fd_sc_hd__a2bb2oi_4 _27380_ (.A1_N(_14329_),
    .A2_N(_10517_),
    .B1(_10514_),
    .B2(_10518_),
    .Y(_10710_));
 sky130_fd_sc_hd__and2_2 _27381_ (.A(_08673_),
    .B(_08085_),
    .X(_10711_));
 sky130_fd_sc_hd__nand3_4 _27382_ (.A(_10515_),
    .B(_09723_),
    .C(_08701_),
    .Y(_10712_));
 sky130_fd_sc_hd__a22o_2 _27383_ (.A1(_07247_),
    .A2(_06940_),
    .B1(_09723_),
    .B2(_07027_),
    .X(_10713_));
 sky130_fd_sc_hd__o21ai_4 _27384_ (.A1(_08699_),
    .A2(_10712_),
    .B1(_10713_),
    .Y(_10714_));
 sky130_fd_sc_hd__xor2_4 _27385_ (.A(_10711_),
    .B(_10714_),
    .X(_10715_));
 sky130_fd_sc_hd__xnor2_4 _27386_ (.A(_10710_),
    .B(_10715_),
    .Y(_10716_));
 sky130_fd_sc_hd__xor2_4 _27387_ (.A(_10709_),
    .B(_10716_),
    .X(_10717_));
 sky130_fd_sc_hd__xnor2_4 _27388_ (.A(_10703_),
    .B(_10717_),
    .Y(_10718_));
 sky130_fd_sc_hd__xor2_4 _27389_ (.A(_10701_),
    .B(_10718_),
    .X(_10719_));
 sky130_fd_sc_hd__o21bai_4 _27390_ (.A1(_10697_),
    .A2(_10699_),
    .B1_N(_10719_),
    .Y(_10720_));
 sky130_fd_sc_hd__nand3b_4 _27391_ (.A_N(_10697_),
    .B(_10719_),
    .C(_10698_),
    .Y(_10721_));
 sky130_fd_sc_hd__nand2_1 _27392_ (.A(_10555_),
    .B(_10528_),
    .Y(_10722_));
 sky130_fd_sc_hd__nand2_4 _27393_ (.A(_10558_),
    .B(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__a21o_1 _27394_ (.A1(_10720_),
    .A2(_10721_),
    .B1(_10723_),
    .X(_10724_));
 sky130_fd_sc_hd__nand3_4 _27395_ (.A(_10723_),
    .B(_10720_),
    .C(_10721_),
    .Y(_10725_));
 sky130_fd_sc_hd__or2b_1 _27396_ (.A(_10586_),
    .B_N(_10574_),
    .X(_10726_));
 sky130_fd_sc_hd__a21boi_4 _27397_ (.A1(_10585_),
    .A2(_10576_),
    .B1_N(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__o22ai_4 _27398_ (.A1(_14276_),
    .A2(_10569_),
    .B1(_10568_),
    .B2(_10571_),
    .Y(_10728_));
 sky130_fd_sc_hd__nand2_1 _27399_ (.A(_07655_),
    .B(_08170_),
    .Y(_10729_));
 sky130_fd_sc_hd__nand3b_4 _27400_ (.A_N(_10729_),
    .B(_12778_),
    .C(_14043_),
    .Y(_10730_));
 sky130_fd_sc_hd__nand2_1 _27401_ (.A(_12777_),
    .B(_09071_),
    .Y(_10731_));
 sky130_fd_sc_hd__nand2_2 _27402_ (.A(_10729_),
    .B(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__nand2_2 _27403_ (.A(_10730_),
    .B(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__xor2_4 _27404_ (.A(_10568_),
    .B(_10733_),
    .X(_10734_));
 sky130_fd_sc_hd__xnor2_4 _27405_ (.A(_10728_),
    .B(_10734_),
    .Y(_10735_));
 sky130_fd_sc_hd__xor2_4 _27406_ (.A(_10415_),
    .B(_10735_),
    .X(_10736_));
 sky130_fd_sc_hd__nor2_1 _27407_ (.A(_10578_),
    .B(_10583_),
    .Y(_10737_));
 sky130_fd_sc_hd__o21bai_4 _27408_ (.A1(_10577_),
    .A2(_10584_),
    .B1_N(_10737_),
    .Y(_10738_));
 sky130_fd_sc_hd__a2bb2oi_4 _27409_ (.A1_N(_14293_),
    .A2_N(_10580_),
    .B1(_10579_),
    .B2(_10581_),
    .Y(_10739_));
 sky130_fd_sc_hd__a2bb2oi_4 _27410_ (.A1_N(_14310_),
    .A2_N(_10509_),
    .B1(_10508_),
    .B2(_10510_),
    .Y(_10740_));
 sky130_fd_sc_hd__and2_2 _27411_ (.A(_05939_),
    .B(_08806_),
    .X(_10741_));
 sky130_fd_sc_hd__nand3_4 _27412_ (.A(_07294_),
    .B(_08721_),
    .C(_07585_),
    .Y(_10742_));
 sky130_fd_sc_hd__a22o_2 _27413_ (.A1(_07294_),
    .A2(_08779_),
    .B1(_08721_),
    .B2(_08487_),
    .X(_10743_));
 sky130_fd_sc_hd__o21ai_4 _27414_ (.A1(_08084_),
    .A2(_10742_),
    .B1(_10743_),
    .Y(_10744_));
 sky130_fd_sc_hd__xor2_4 _27415_ (.A(_10741_),
    .B(_10744_),
    .X(_10745_));
 sky130_fd_sc_hd__xnor2_4 _27416_ (.A(_10740_),
    .B(_10745_),
    .Y(_10746_));
 sky130_fd_sc_hd__xor2_4 _27417_ (.A(_10739_),
    .B(_10746_),
    .X(_10747_));
 sky130_fd_sc_hd__xnor2_4 _27418_ (.A(_10738_),
    .B(_10747_),
    .Y(_10748_));
 sky130_fd_sc_hd__xnor2_4 _27419_ (.A(_10736_),
    .B(_10748_),
    .Y(_10749_));
 sky130_fd_sc_hd__and2_1 _27420_ (.A(_10524_),
    .B(_10522_),
    .X(_10750_));
 sky130_fd_sc_hd__o21bai_4 _27421_ (.A1(_10507_),
    .A2(_10525_),
    .B1_N(_10750_),
    .Y(_10751_));
 sky130_fd_sc_hd__xnor2_4 _27422_ (.A(_10749_),
    .B(_10751_),
    .Y(_10752_));
 sky130_fd_sc_hd__xnor2_4 _27423_ (.A(_10727_),
    .B(_10752_),
    .Y(_10753_));
 sky130_fd_sc_hd__a21boi_2 _27424_ (.A1(_10724_),
    .A2(_10725_),
    .B1_N(_10753_),
    .Y(_10754_));
 sky130_fd_sc_hd__nand3b_4 _27425_ (.A_N(_10753_),
    .B(_10724_),
    .C(_10725_),
    .Y(_10755_));
 sky130_vsdinv _27426_ (.A(_10755_),
    .Y(_10756_));
 sky130_fd_sc_hd__nand2_4 _27427_ (.A(_10595_),
    .B(_10561_),
    .Y(_10757_));
 sky130_fd_sc_hd__o21bai_4 _27428_ (.A1(_10754_),
    .A2(_10756_),
    .B1_N(_10757_),
    .Y(_10758_));
 sky130_fd_sc_hd__a21bo_1 _27429_ (.A1(_10724_),
    .A2(_10725_),
    .B1_N(_10753_),
    .X(_10759_));
 sky130_fd_sc_hd__nand3_4 _27430_ (.A(_10757_),
    .B(_10759_),
    .C(_10755_),
    .Y(_10760_));
 sky130_vsdinv _27431_ (.A(_10590_),
    .Y(_10761_));
 sky130_fd_sc_hd__nor2_2 _27432_ (.A(_10606_),
    .B(_10613_),
    .Y(_10762_));
 sky130_fd_sc_hd__a21oi_4 _27433_ (.A1(_10608_),
    .A2(_10612_),
    .B1(_10762_),
    .Y(_10763_));
 sky130_fd_sc_hd__or2_4 _27434_ (.A(_10610_),
    .B(_09968_),
    .X(_10764_));
 sky130_fd_sc_hd__and2_1 _27435_ (.A(_09968_),
    .B(_10610_),
    .X(_10765_));
 sky130_fd_sc_hd__a21oi_4 _27436_ (.A1(_10764_),
    .A2(_10609_),
    .B1(_10765_),
    .Y(_10766_));
 sky130_fd_sc_hd__nor2_1 _27437_ (.A(_10567_),
    .B(_10572_),
    .Y(_10767_));
 sky130_fd_sc_hd__o21bai_4 _27438_ (.A1(_10415_),
    .A2(_10573_),
    .B1_N(_10767_),
    .Y(_10768_));
 sky130_fd_sc_hd__xnor2_4 _27439_ (.A(_10768_),
    .B(_10612_),
    .Y(_10769_));
 sky130_fd_sc_hd__xor2_4 _27440_ (.A(_10766_),
    .B(_10769_),
    .X(_10770_));
 sky130_fd_sc_hd__xor2_4 _27441_ (.A(_10763_),
    .B(_10770_),
    .X(_10771_));
 sky130_fd_sc_hd__nor2_2 _27442_ (.A(_10149_),
    .B(_10771_),
    .Y(_10772_));
 sky130_fd_sc_hd__and2_1 _27443_ (.A(_10771_),
    .B(_09793_),
    .X(_10773_));
 sky130_fd_sc_hd__a211o_1 _27444_ (.A1(_10761_),
    .A2(_10589_),
    .B1(_10772_),
    .C1(_10773_),
    .X(_10774_));
 sky130_fd_sc_hd__o211ai_4 _27445_ (.A1(_10772_),
    .A2(_10773_),
    .B1(_10589_),
    .C1(_10761_),
    .Y(_10775_));
 sky130_fd_sc_hd__or2b_1 _27446_ (.A(_10604_),
    .B_N(_10614_),
    .X(_10776_));
 sky130_fd_sc_hd__o21a_1 _27447_ (.A1(_10149_),
    .A2(_10615_),
    .B1(_10776_),
    .X(_10777_));
 sky130_vsdinv _27448_ (.A(_10777_),
    .Y(_10778_));
 sky130_fd_sc_hd__a21oi_4 _27449_ (.A1(_10774_),
    .A2(_10775_),
    .B1(_10778_),
    .Y(_10779_));
 sky130_fd_sc_hd__and3_1 _27450_ (.A(_10774_),
    .B(_10775_),
    .C(_10778_),
    .X(_10780_));
 sky130_fd_sc_hd__nor2_4 _27451_ (.A(_10779_),
    .B(_10780_),
    .Y(_10781_));
 sky130_fd_sc_hd__a21oi_2 _27452_ (.A1(_10758_),
    .A2(_10760_),
    .B1(_10781_),
    .Y(_10782_));
 sky130_vsdinv _27453_ (.A(_10781_),
    .Y(_10783_));
 sky130_fd_sc_hd__a21oi_4 _27454_ (.A1(_10759_),
    .A2(_10755_),
    .B1(_10757_),
    .Y(_10784_));
 sky130_fd_sc_hd__nor3b_4 _27455_ (.A(_10783_),
    .B(_10784_),
    .C_N(_10760_),
    .Y(_10785_));
 sky130_vsdinv _27456_ (.A(_10625_),
    .Y(_10786_));
 sky130_fd_sc_hd__a21oi_4 _27457_ (.A1(_10599_),
    .A2(_10595_),
    .B1(_10597_),
    .Y(_10787_));
 sky130_fd_sc_hd__o21ai_4 _27458_ (.A1(_10786_),
    .A2(_10787_),
    .B1(_10600_),
    .Y(_10788_));
 sky130_fd_sc_hd__o21bai_4 _27459_ (.A1(_10782_),
    .A2(_10785_),
    .B1_N(_10788_),
    .Y(_10789_));
 sky130_fd_sc_hd__o2bb2ai_2 _27460_ (.A1_N(_10760_),
    .A2_N(_10758_),
    .B1(_10780_),
    .B2(_10779_),
    .Y(_10790_));
 sky130_fd_sc_hd__nand3_4 _27461_ (.A(_10758_),
    .B(_10781_),
    .C(_10760_),
    .Y(_10791_));
 sky130_fd_sc_hd__nand3_4 _27462_ (.A(_10790_),
    .B(_10791_),
    .C(_10788_),
    .Y(_10792_));
 sky130_fd_sc_hd__o21ai_4 _27463_ (.A1(_10602_),
    .A2(_10624_),
    .B1(_10622_),
    .Y(_10793_));
 sky130_fd_sc_hd__xor2_4 _27464_ (.A(net414),
    .B(_10793_),
    .X(_10794_));
 sky130_fd_sc_hd__a21oi_2 _27465_ (.A1(_10789_),
    .A2(_10792_),
    .B1(_10794_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand3_4 _27466_ (.A(_10789_),
    .B(_10794_),
    .C(_10792_),
    .Y(_10796_));
 sky130_vsdinv _27467_ (.A(_10796_),
    .Y(_10797_));
 sky130_vsdinv _27468_ (.A(_10637_),
    .Y(_10798_));
 sky130_fd_sc_hd__a21oi_1 _27469_ (.A1(_10626_),
    .A2(_10627_),
    .B1(_10628_),
    .Y(_10799_));
 sky130_fd_sc_hd__o21ai_2 _27470_ (.A1(_10798_),
    .A2(_10799_),
    .B1(_10629_),
    .Y(_10800_));
 sky130_fd_sc_hd__o21bai_4 _27471_ (.A1(_10795_),
    .A2(_10797_),
    .B1_N(_10800_),
    .Y(_10801_));
 sky130_fd_sc_hd__and2_1 _27472_ (.A(_10793_),
    .B(net414),
    .X(_10802_));
 sky130_fd_sc_hd__o211a_1 _27473_ (.A1(_10602_),
    .A2(_10624_),
    .B1(_10325_),
    .C1(_10622_),
    .X(_10803_));
 sky130_fd_sc_hd__o2bb2ai_2 _27474_ (.A1_N(_10792_),
    .A2_N(_10789_),
    .B1(_10802_),
    .B2(_10803_),
    .Y(_10804_));
 sky130_fd_sc_hd__nand3_4 _27475_ (.A(_10804_),
    .B(_10796_),
    .C(_10800_),
    .Y(_10805_));
 sky130_fd_sc_hd__a21oi_2 _27476_ (.A1(_10801_),
    .A2(_10805_),
    .B1(_10634_),
    .Y(_10806_));
 sky130_fd_sc_hd__nand3_4 _27477_ (.A(_10801_),
    .B(_10634_),
    .C(_10805_),
    .Y(_10807_));
 sky130_vsdinv _27478_ (.A(_10807_),
    .Y(_10808_));
 sky130_vsdinv _27479_ (.A(_10643_),
    .Y(_10809_));
 sky130_fd_sc_hd__o21ai_4 _27480_ (.A1(_10809_),
    .A2(_10640_),
    .B1(_10641_),
    .Y(_10810_));
 sky130_fd_sc_hd__o21bai_1 _27481_ (.A1(_10806_),
    .A2(_10808_),
    .B1_N(_10810_),
    .Y(_10811_));
 sky130_fd_sc_hd__buf_6 _27482_ (.A(_10338_),
    .X(_10812_));
 sky130_fd_sc_hd__buf_6 _27483_ (.A(_10812_),
    .X(_10813_));
 sky130_fd_sc_hd__o2bb2ai_4 _27484_ (.A1_N(_10805_),
    .A2_N(_10801_),
    .B1(_10813_),
    .B2(_10633_),
    .Y(_10814_));
 sky130_fd_sc_hd__nand3_4 _27485_ (.A(_10814_),
    .B(_10810_),
    .C(_10807_),
    .Y(_10815_));
 sky130_fd_sc_hd__nand2_1 _27486_ (.A(_10811_),
    .B(_10815_),
    .Y(_10816_));
 sky130_fd_sc_hd__a21oi_1 _27487_ (.A1(_10647_),
    .A2(_10641_),
    .B1(_10643_),
    .Y(_10817_));
 sky130_vsdinv _27488_ (.A(_10648_),
    .Y(_10818_));
 sky130_fd_sc_hd__o21bai_1 _27489_ (.A1(_10817_),
    .A2(_10818_),
    .B1_N(_10650_),
    .Y(_10819_));
 sky130_fd_sc_hd__a21oi_1 _27490_ (.A1(_10666_),
    .A2(_10819_),
    .B1(_10653_),
    .Y(_10820_));
 sky130_fd_sc_hd__xor2_1 _27491_ (.A(_10816_),
    .B(_10820_),
    .X(_02664_));
 sky130_fd_sc_hd__nor2_1 _27492_ (.A(_10710_),
    .B(_10715_),
    .Y(_10821_));
 sky130_fd_sc_hd__o21ba_1 _27493_ (.A1(_10709_),
    .A2(_10716_),
    .B1_N(_10821_),
    .X(_10822_));
 sky130_fd_sc_hd__nor2_1 _27494_ (.A(_10670_),
    .B(_10676_),
    .Y(_10823_));
 sky130_fd_sc_hd__o21bai_4 _27495_ (.A1(_10669_),
    .A2(_10677_),
    .B1_N(_10823_),
    .Y(_10824_));
 sky130_fd_sc_hd__buf_2 _27496_ (.A(_07778_),
    .X(_10825_));
 sky130_fd_sc_hd__and2_2 _27497_ (.A(_06061_),
    .B(_10825_),
    .X(_10826_));
 sky130_fd_sc_hd__clkbuf_4 _27498_ (.A(_07477_),
    .X(_10827_));
 sky130_fd_sc_hd__nand3_4 _27499_ (.A(_08857_),
    .B(_10705_),
    .C(_10827_),
    .Y(_10828_));
 sky130_fd_sc_hd__buf_2 _27500_ (.A(_07578_),
    .X(_10829_));
 sky130_fd_sc_hd__a22o_2 _27501_ (.A1(_08857_),
    .A2(_10827_),
    .B1(_08423_),
    .B2(_10829_),
    .X(_10830_));
 sky130_fd_sc_hd__o21ai_4 _27502_ (.A1(_14298_),
    .A2(_10828_),
    .B1(_10830_),
    .Y(_10831_));
 sky130_fd_sc_hd__xor2_4 _27503_ (.A(_10826_),
    .B(_10831_),
    .X(_10832_));
 sky130_fd_sc_hd__a2bb2oi_4 _27504_ (.A1_N(_14321_),
    .A2_N(_10712_),
    .B1(_10711_),
    .B2(_10713_),
    .Y(_10833_));
 sky130_fd_sc_hd__and2_2 _27505_ (.A(_06471_),
    .B(_07210_),
    .X(_10834_));
 sky130_fd_sc_hd__nand3_4 _27506_ (.A(_07247_),
    .B(_09723_),
    .C(_07027_),
    .Y(_10835_));
 sky130_fd_sc_hd__a22o_2 _27507_ (.A1(_09197_),
    .A2(_07036_),
    .B1(_08668_),
    .B2(_07039_),
    .X(_10836_));
 sky130_fd_sc_hd__o21ai_4 _27508_ (.A1(_14314_),
    .A2(_10835_),
    .B1(_10836_),
    .Y(_10837_));
 sky130_fd_sc_hd__xor2_4 _27509_ (.A(_10834_),
    .B(_10837_),
    .X(_10838_));
 sky130_fd_sc_hd__xnor2_4 _27510_ (.A(_10833_),
    .B(_10838_),
    .Y(_10839_));
 sky130_fd_sc_hd__xor2_4 _27511_ (.A(_10832_),
    .B(_10839_),
    .X(_10840_));
 sky130_fd_sc_hd__xnor2_2 _27512_ (.A(_10824_),
    .B(_10840_),
    .Y(_10841_));
 sky130_fd_sc_hd__xor2_2 _27513_ (.A(_10822_),
    .B(_10841_),
    .X(_10842_));
 sky130_vsdinv _27514_ (.A(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__and2_1 _27515_ (.A(_10694_),
    .B(_10680_),
    .X(_10844_));
 sky130_fd_sc_hd__o21bai_2 _27516_ (.A1(_10678_),
    .A2(_10695_),
    .B1_N(_10844_),
    .Y(_10845_));
 sky130_fd_sc_hd__a2bb2oi_4 _27517_ (.A1_N(_14342_),
    .A2_N(_10673_),
    .B1(_10671_),
    .B2(_10674_),
    .Y(_10846_));
 sky130_fd_sc_hd__a2bb2oi_4 _27518_ (.A1_N(_14361_),
    .A2_N(_10682_),
    .B1(_10681_),
    .B2(_10683_),
    .Y(_10847_));
 sky130_fd_sc_hd__and2_2 _27519_ (.A(_06888_),
    .B(_07034_),
    .X(_10848_));
 sky130_fd_sc_hd__nand3_4 _27520_ (.A(_10672_),
    .B(_07103_),
    .C(_07747_),
    .Y(_10849_));
 sky130_fd_sc_hd__a22o_2 _27521_ (.A1(_09152_),
    .A2(_06441_),
    .B1(_09153_),
    .B2(_06761_),
    .X(_10850_));
 sky130_fd_sc_hd__o21ai_4 _27522_ (.A1(_07214_),
    .A2(_10849_),
    .B1(_10850_),
    .Y(_10851_));
 sky130_fd_sc_hd__xor2_4 _27523_ (.A(_10848_),
    .B(_10851_),
    .X(_10852_));
 sky130_fd_sc_hd__xnor2_4 _27524_ (.A(_10847_),
    .B(_10852_),
    .Y(_10853_));
 sky130_fd_sc_hd__xnor2_4 _27525_ (.A(_10846_),
    .B(_10853_),
    .Y(_10854_));
 sky130_fd_sc_hd__or2b_1 _27526_ (.A(_10692_),
    .B_N(_10687_),
    .X(_10855_));
 sky130_fd_sc_hd__o21ai_4 _27527_ (.A1(_10685_),
    .A2(_10693_),
    .B1(_10855_),
    .Y(_10856_));
 sky130_fd_sc_hd__and2_2 _27528_ (.A(_07873_),
    .B(_06432_),
    .X(_10857_));
 sky130_fd_sc_hd__nand3_4 _27529_ (.A(_13972_),
    .B(_13978_),
    .C(_06147_),
    .Y(_10858_));
 sky130_fd_sc_hd__a22o_2 _27530_ (.A1(_09357_),
    .A2(_06030_),
    .B1(_09162_),
    .B2(_06279_),
    .X(_10859_));
 sky130_fd_sc_hd__o21ai_4 _27531_ (.A1(_08338_),
    .A2(_10858_),
    .B1(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__xor2_4 _27532_ (.A(_10857_),
    .B(_10860_),
    .X(_10861_));
 sky130_fd_sc_hd__nand3b_4 _27533_ (.A_N(_10689_),
    .B(_09876_),
    .C(_14384_),
    .Y(_10862_));
 sky130_fd_sc_hd__o31ai_4 _27534_ (.A1(_13967_),
    .A2(_14373_),
    .A3(_10691_),
    .B1(_10862_),
    .Y(_10863_));
 sky130_fd_sc_hd__and2_2 _27535_ (.A(_07945_),
    .B(_08720_),
    .X(_10864_));
 sky130_fd_sc_hd__nand2_2 _27536_ (.A(_13961_),
    .B(_05768_),
    .Y(_10865_));
 sky130_fd_sc_hd__and2b_1 _27537_ (.A_N(_05690_),
    .B(_12804_),
    .X(_10866_));
 sky130_fd_sc_hd__xor2_4 _27538_ (.A(_10865_),
    .B(_10866_),
    .X(_10867_));
 sky130_fd_sc_hd__xor2_4 _27539_ (.A(_10864_),
    .B(_10867_),
    .X(_10868_));
 sky130_fd_sc_hd__xor2_4 _27540_ (.A(_10863_),
    .B(_10868_),
    .X(_10869_));
 sky130_fd_sc_hd__xor2_4 _27541_ (.A(_10861_),
    .B(_10869_),
    .X(_10870_));
 sky130_fd_sc_hd__xnor2_4 _27542_ (.A(_10856_),
    .B(_10870_),
    .Y(_10871_));
 sky130_fd_sc_hd__xor2_4 _27543_ (.A(_10854_),
    .B(_10871_),
    .X(_10872_));
 sky130_fd_sc_hd__xnor2_1 _27544_ (.A(_10845_),
    .B(_10872_),
    .Y(_10873_));
 sky130_fd_sc_hd__nor2_2 _27545_ (.A(_10843_),
    .B(_10873_),
    .Y(_10874_));
 sky130_fd_sc_hd__and2_1 _27546_ (.A(_10873_),
    .B(_10843_),
    .X(_10875_));
 sky130_fd_sc_hd__nand2_1 _27547_ (.A(_10721_),
    .B(_10698_),
    .Y(_10876_));
 sky130_fd_sc_hd__o21ba_1 _27548_ (.A1(_10874_),
    .A2(_10875_),
    .B1_N(_10876_),
    .X(_10877_));
 sky130_vsdinv _27549_ (.A(_10877_),
    .Y(_10878_));
 sky130_fd_sc_hd__a211o_4 _27550_ (.A1(_10698_),
    .A2(_10721_),
    .B1(_10874_),
    .C1(_10875_),
    .X(_10879_));
 sky130_fd_sc_hd__and2b_1 _27551_ (.A_N(_10748_),
    .B(_10736_),
    .X(_10880_));
 sky130_fd_sc_hd__a21oi_4 _27552_ (.A1(_10747_),
    .A2(_10738_),
    .B1(_10880_),
    .Y(_10881_));
 sky130_fd_sc_hd__and2_1 _27553_ (.A(_10717_),
    .B(_10703_),
    .X(_10882_));
 sky130_fd_sc_hd__o21bai_4 _27554_ (.A1(_10701_),
    .A2(_10718_),
    .B1_N(_10882_),
    .Y(_10883_));
 sky130_fd_sc_hd__o21ai_2 _27555_ (.A1(_14038_),
    .A2(_14043_),
    .B1(_09468_),
    .Y(_10884_));
 sky130_fd_sc_hd__nand3_4 _27556_ (.A(_09468_),
    .B(_14038_),
    .C(_14043_),
    .Y(_10885_));
 sky130_fd_sc_hd__and2b_2 _27557_ (.A_N(_10884_),
    .B(_10885_),
    .X(_10886_));
 sky130_fd_sc_hd__a22oi_4 _27558_ (.A1(_05442_),
    .A2(_10732_),
    .B1(_10730_),
    .B2(_10568_),
    .Y(_10887_));
 sky130_fd_sc_hd__xor2_4 _27559_ (.A(_10886_),
    .B(_10887_),
    .X(_10888_));
 sky130_fd_sc_hd__xor2_4 _27560_ (.A(_10414_),
    .B(_10888_),
    .X(_10889_));
 sky130_fd_sc_hd__nor2_1 _27561_ (.A(_10740_),
    .B(_10745_),
    .Y(_10890_));
 sky130_fd_sc_hd__o21bai_4 _27562_ (.A1(_10739_),
    .A2(_10746_),
    .B1_N(_10890_),
    .Y(_10891_));
 sky130_fd_sc_hd__a2bb2oi_4 _27563_ (.A1_N(_14287_),
    .A2_N(_10742_),
    .B1(_10741_),
    .B2(_10743_),
    .Y(_10892_));
 sky130_fd_sc_hd__a2bb2oi_4 _27564_ (.A1_N(_09222_),
    .A2_N(_10706_),
    .B1(_10704_),
    .B2(_10707_),
    .Y(_10893_));
 sky130_fd_sc_hd__and2_2 _27565_ (.A(_05939_),
    .B(_08595_),
    .X(_10894_));
 sky130_fd_sc_hd__nand3_4 _27566_ (.A(_07820_),
    .B(_08721_),
    .C(_08073_),
    .Y(_10895_));
 sky130_fd_sc_hd__a22o_2 _27567_ (.A1(_07294_),
    .A2(_08487_),
    .B1(_08721_),
    .B2(_08165_),
    .X(_10896_));
 sky130_fd_sc_hd__o21ai_4 _27568_ (.A1(_14279_),
    .A2(_10895_),
    .B1(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__xor2_4 _27569_ (.A(_10894_),
    .B(_10897_),
    .X(_10898_));
 sky130_fd_sc_hd__xnor2_4 _27570_ (.A(_10893_),
    .B(_10898_),
    .Y(_10899_));
 sky130_fd_sc_hd__xor2_4 _27571_ (.A(_10892_),
    .B(_10899_),
    .X(_10900_));
 sky130_fd_sc_hd__xnor2_4 _27572_ (.A(_10891_),
    .B(_10900_),
    .Y(_10901_));
 sky130_fd_sc_hd__xnor2_4 _27573_ (.A(_10889_),
    .B(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__xnor2_2 _27574_ (.A(_10883_),
    .B(_10902_),
    .Y(_10903_));
 sky130_fd_sc_hd__xnor2_2 _27575_ (.A(_10881_),
    .B(_10903_),
    .Y(_10904_));
 sky130_fd_sc_hd__a21boi_2 _27576_ (.A1(_10878_),
    .A2(_10879_),
    .B1_N(_10904_),
    .Y(_10905_));
 sky130_fd_sc_hd__nand3b_4 _27577_ (.A_N(_10904_),
    .B(_10878_),
    .C(_10879_),
    .Y(_10906_));
 sky130_vsdinv _27578_ (.A(_10906_),
    .Y(_10907_));
 sky130_fd_sc_hd__a21oi_2 _27579_ (.A1(_10720_),
    .A2(_10721_),
    .B1(_10723_),
    .Y(_10908_));
 sky130_fd_sc_hd__o21ai_4 _27580_ (.A1(_10753_),
    .A2(_10908_),
    .B1(_10725_),
    .Y(_10909_));
 sky130_fd_sc_hd__o21bai_4 _27581_ (.A1(_10905_),
    .A2(_10907_),
    .B1_N(_10909_),
    .Y(_10910_));
 sky130_fd_sc_hd__a21bo_2 _27582_ (.A1(_10878_),
    .A2(_10879_),
    .B1_N(_10904_),
    .X(_10911_));
 sky130_fd_sc_hd__nand3_4 _27583_ (.A(_10911_),
    .B(_10906_),
    .C(_10909_),
    .Y(_10912_));
 sky130_vsdinv _27584_ (.A(_10766_),
    .Y(_10913_));
 sky130_fd_sc_hd__and2_1 _27585_ (.A(_10734_),
    .B(_10728_),
    .X(_10914_));
 sky130_fd_sc_hd__o21bai_4 _27586_ (.A1(_10415_),
    .A2(_10735_),
    .B1_N(_10914_),
    .Y(_10915_));
 sky130_fd_sc_hd__xor2_4 _27587_ (.A(_10915_),
    .B(_10612_),
    .X(_10916_));
 sky130_fd_sc_hd__xor2_4 _27588_ (.A(_10913_),
    .B(_10916_),
    .X(_10917_));
 sky130_fd_sc_hd__nor2_1 _27589_ (.A(_10766_),
    .B(_10769_),
    .Y(_10918_));
 sky130_fd_sc_hd__a21o_1 _27590_ (.A1(_10612_),
    .A2(_10768_),
    .B1(_10918_),
    .X(_10919_));
 sky130_fd_sc_hd__nor2_4 _27591_ (.A(_10917_),
    .B(_10919_),
    .Y(_10920_));
 sky130_fd_sc_hd__and2_1 _27592_ (.A(_10919_),
    .B(_10917_),
    .X(_10921_));
 sky130_fd_sc_hd__nor3_4 _27593_ (.A(_10446_),
    .B(_10920_),
    .C(_10921_),
    .Y(_10922_));
 sky130_fd_sc_hd__o21a_1 _27594_ (.A1(_10920_),
    .A2(_10921_),
    .B1(_09985_),
    .X(_10923_));
 sky130_fd_sc_hd__nand2_1 _27595_ (.A(_10751_),
    .B(_10749_),
    .Y(_10924_));
 sky130_fd_sc_hd__o21a_1 _27596_ (.A1(_10727_),
    .A2(_10752_),
    .B1(_10924_),
    .X(_10925_));
 sky130_fd_sc_hd__or3_4 _27597_ (.A(_10922_),
    .B(_10923_),
    .C(_10925_),
    .X(_10926_));
 sky130_fd_sc_hd__o21ai_4 _27598_ (.A1(_10922_),
    .A2(_10923_),
    .B1(_10925_),
    .Y(_10927_));
 sky130_fd_sc_hd__and2b_1 _27599_ (.A_N(_10763_),
    .B(_10770_),
    .X(_10928_));
 sky130_fd_sc_hd__o21ba_1 _27600_ (.A1(_10446_),
    .A2(_10771_),
    .B1_N(_10928_),
    .X(_10929_));
 sky130_vsdinv _27601_ (.A(_10929_),
    .Y(_10930_));
 sky130_fd_sc_hd__a21oi_1 _27602_ (.A1(_10926_),
    .A2(_10927_),
    .B1(_10930_),
    .Y(_10931_));
 sky130_fd_sc_hd__nand3_4 _27603_ (.A(_10926_),
    .B(_10930_),
    .C(_10927_),
    .Y(_10932_));
 sky130_fd_sc_hd__and2b_1 _27604_ (.A_N(_10931_),
    .B(_10932_),
    .X(_10933_));
 sky130_fd_sc_hd__a21oi_2 _27605_ (.A1(_10910_),
    .A2(_10912_),
    .B1(_10933_),
    .Y(_10934_));
 sky130_fd_sc_hd__or2b_2 _27606_ (.A(_10931_),
    .B_N(_10932_),
    .X(_10935_));
 sky130_fd_sc_hd__a21oi_4 _27607_ (.A1(_10911_),
    .A2(_10906_),
    .B1(_10909_),
    .Y(_10936_));
 sky130_vsdinv _27608_ (.A(_10912_),
    .Y(_10937_));
 sky130_fd_sc_hd__nor3_4 _27609_ (.A(_10935_),
    .B(_10936_),
    .C(_10937_),
    .Y(_10938_));
 sky130_fd_sc_hd__o21ai_4 _27610_ (.A1(_10783_),
    .A2(_10784_),
    .B1(_10760_),
    .Y(_10939_));
 sky130_fd_sc_hd__o21bai_4 _27611_ (.A1(_10934_),
    .A2(_10938_),
    .B1_N(_10939_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand2_1 _27612_ (.A(_10910_),
    .B(_10912_),
    .Y(_10941_));
 sky130_fd_sc_hd__nand2_2 _27613_ (.A(_10941_),
    .B(_10935_),
    .Y(_10942_));
 sky130_fd_sc_hd__nand3_4 _27614_ (.A(_10910_),
    .B(_10933_),
    .C(_10912_),
    .Y(_10943_));
 sky130_fd_sc_hd__nand3_4 _27615_ (.A(_10942_),
    .B(_10943_),
    .C(_10939_),
    .Y(_10944_));
 sky130_fd_sc_hd__a21bo_2 _27616_ (.A1(_10778_),
    .A2(_10775_),
    .B1_N(_10774_),
    .X(_10945_));
 sky130_fd_sc_hd__xor2_4 _27617_ (.A(net414),
    .B(_10945_),
    .X(_10946_));
 sky130_fd_sc_hd__a21oi_4 _27618_ (.A1(_10940_),
    .A2(_10944_),
    .B1(_10946_),
    .Y(_10947_));
 sky130_vsdinv _27619_ (.A(_10946_),
    .Y(_10948_));
 sky130_fd_sc_hd__a21oi_4 _27620_ (.A1(_10942_),
    .A2(_10943_),
    .B1(_10939_),
    .Y(_10949_));
 sky130_vsdinv _27621_ (.A(_10944_),
    .Y(_10950_));
 sky130_fd_sc_hd__nor3_4 _27622_ (.A(_10948_),
    .B(_10949_),
    .C(_10950_),
    .Y(_10951_));
 sky130_vsdinv _27623_ (.A(_10794_),
    .Y(_10952_));
 sky130_fd_sc_hd__a21oi_2 _27624_ (.A1(_10790_),
    .A2(_10791_),
    .B1(_10788_),
    .Y(_10953_));
 sky130_fd_sc_hd__o21ai_4 _27625_ (.A1(_10952_),
    .A2(_10953_),
    .B1(_10792_),
    .Y(_10954_));
 sky130_fd_sc_hd__o21bai_1 _27626_ (.A1(_10947_),
    .A2(_10951_),
    .B1_N(_10954_),
    .Y(_10955_));
 sky130_fd_sc_hd__nand2_1 _27627_ (.A(_10940_),
    .B(_10944_),
    .Y(_10956_));
 sky130_fd_sc_hd__nand2_2 _27628_ (.A(_10956_),
    .B(_10948_),
    .Y(_10957_));
 sky130_fd_sc_hd__nand3_4 _27629_ (.A(_10940_),
    .B(_10946_),
    .C(_10944_),
    .Y(_10958_));
 sky130_fd_sc_hd__nand3_2 _27630_ (.A(_10957_),
    .B(_10954_),
    .C(_10958_),
    .Y(_10959_));
 sky130_fd_sc_hd__a21oi_1 _27631_ (.A1(_10955_),
    .A2(_10959_),
    .B1(_10802_),
    .Y(_10960_));
 sky130_vsdinv _27632_ (.A(_10802_),
    .Y(_10961_));
 sky130_fd_sc_hd__a21oi_4 _27633_ (.A1(_10957_),
    .A2(_10958_),
    .B1(_10954_),
    .Y(_10962_));
 sky130_fd_sc_hd__a21boi_4 _27634_ (.A1(_10789_),
    .A2(_10794_),
    .B1_N(_10792_),
    .Y(_10963_));
 sky130_fd_sc_hd__nor3_4 _27635_ (.A(_10947_),
    .B(_10963_),
    .C(_10951_),
    .Y(_10964_));
 sky130_fd_sc_hd__nor3_2 _27636_ (.A(_10961_),
    .B(_10962_),
    .C(_10964_),
    .Y(_10965_));
 sky130_vsdinv _27637_ (.A(_10634_),
    .Y(_10966_));
 sky130_fd_sc_hd__a21oi_1 _27638_ (.A1(_10804_),
    .A2(_10796_),
    .B1(_10800_),
    .Y(_10967_));
 sky130_fd_sc_hd__o21ai_1 _27639_ (.A1(_10966_),
    .A2(_10967_),
    .B1(_10805_),
    .Y(_10968_));
 sky130_fd_sc_hd__o21bai_1 _27640_ (.A1(_10960_),
    .A2(_10965_),
    .B1_N(_10968_),
    .Y(_10969_));
 sky130_fd_sc_hd__o21bai_1 _27641_ (.A1(_10962_),
    .A2(_10964_),
    .B1_N(_10802_),
    .Y(_10970_));
 sky130_fd_sc_hd__nand3_1 _27642_ (.A(_10955_),
    .B(_10802_),
    .C(_10959_),
    .Y(_10971_));
 sky130_fd_sc_hd__nand3_2 _27643_ (.A(_10970_),
    .B(_10968_),
    .C(_10971_),
    .Y(_10972_));
 sky130_fd_sc_hd__nand2_1 _27644_ (.A(_10969_),
    .B(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__nand2_1 _27645_ (.A(_10819_),
    .B(_10652_),
    .Y(_10974_));
 sky130_fd_sc_hd__nor2_2 _27646_ (.A(_10974_),
    .B(_10816_),
    .Y(_10975_));
 sky130_fd_sc_hd__a21oi_4 _27647_ (.A1(_10814_),
    .A2(_10807_),
    .B1(_10810_),
    .Y(_10976_));
 sky130_fd_sc_hd__a21oi_4 _27648_ (.A1(_10652_),
    .A2(_10815_),
    .B1(_10976_),
    .Y(_10977_));
 sky130_fd_sc_hd__a21oi_2 _27649_ (.A1(_10666_),
    .A2(_10975_),
    .B1(_10977_),
    .Y(_10978_));
 sky130_fd_sc_hd__xor2_1 _27650_ (.A(_10973_),
    .B(_10978_),
    .X(_02665_));
 sky130_fd_sc_hd__nor2_1 _27651_ (.A(_10833_),
    .B(_10838_),
    .Y(_10979_));
 sky130_fd_sc_hd__o21ba_1 _27652_ (.A1(_10832_),
    .A2(_10839_),
    .B1_N(_10979_),
    .X(_10980_));
 sky130_fd_sc_hd__nor2_1 _27653_ (.A(_10847_),
    .B(_10852_),
    .Y(_10981_));
 sky130_fd_sc_hd__o21bai_2 _27654_ (.A1(_10846_),
    .A2(_10853_),
    .B1_N(_10981_),
    .Y(_10982_));
 sky130_fd_sc_hd__and2_2 _27655_ (.A(_06061_),
    .B(_08489_),
    .X(_10983_));
 sky130_fd_sc_hd__buf_2 _27656_ (.A(_08425_),
    .X(_10984_));
 sky130_fd_sc_hd__nand3_4 _27657_ (.A(_10984_),
    .B(_10705_),
    .C(_07770_),
    .Y(_10985_));
 sky130_fd_sc_hd__a22o_2 _27658_ (.A1(_10984_),
    .A2(_07770_),
    .B1(_10705_),
    .B2(_10825_),
    .X(_10986_));
 sky130_fd_sc_hd__o21ai_4 _27659_ (.A1(_14294_),
    .A2(_10985_),
    .B1(_10986_),
    .Y(_10987_));
 sky130_fd_sc_hd__xor2_4 _27660_ (.A(_10983_),
    .B(_10987_),
    .X(_10988_));
 sky130_fd_sc_hd__a2bb2oi_4 _27661_ (.A1_N(_14316_),
    .A2_N(_10835_),
    .B1(_10834_),
    .B2(_10836_),
    .Y(_10989_));
 sky130_fd_sc_hd__and2_2 _27662_ (.A(_06472_),
    .B(_07570_),
    .X(_10990_));
 sky130_fd_sc_hd__buf_4 _27663_ (.A(_09197_),
    .X(_10991_));
 sky130_fd_sc_hd__buf_4 _27664_ (.A(_09723_),
    .X(_10992_));
 sky130_fd_sc_hd__nand3_4 _27665_ (.A(_10991_),
    .B(_10992_),
    .C(_07199_),
    .Y(_10993_));
 sky130_fd_sc_hd__a22o_2 _27666_ (.A1(_10991_),
    .A2(_07473_),
    .B1(_10992_),
    .B2(_07575_),
    .X(_10994_));
 sky130_fd_sc_hd__o21ai_4 _27667_ (.A1(_14310_),
    .A2(_10993_),
    .B1(_10994_),
    .Y(_10995_));
 sky130_fd_sc_hd__xor2_4 _27668_ (.A(_10990_),
    .B(_10995_),
    .X(_10996_));
 sky130_fd_sc_hd__xnor2_4 _27669_ (.A(_10989_),
    .B(_10996_),
    .Y(_10997_));
 sky130_fd_sc_hd__xor2_4 _27670_ (.A(_10988_),
    .B(_10997_),
    .X(_10998_));
 sky130_fd_sc_hd__xnor2_2 _27671_ (.A(_10982_),
    .B(_10998_),
    .Y(_10999_));
 sky130_fd_sc_hd__xor2_1 _27672_ (.A(_10980_),
    .B(_10999_),
    .X(_11000_));
 sky130_fd_sc_hd__and2_1 _27673_ (.A(_10870_),
    .B(_10856_),
    .X(_11001_));
 sky130_fd_sc_hd__o21bai_1 _27674_ (.A1(_10854_),
    .A2(_10871_),
    .B1_N(_11001_),
    .Y(_11002_));
 sky130_fd_sc_hd__a2bb2oi_4 _27675_ (.A1_N(_14335_),
    .A2_N(_10849_),
    .B1(_10848_),
    .B2(_10850_),
    .Y(_11003_));
 sky130_fd_sc_hd__a2bb2oi_4 _27676_ (.A1_N(_14354_),
    .A2_N(_10858_),
    .B1(_10857_),
    .B2(_10859_),
    .Y(_11004_));
 sky130_fd_sc_hd__and2_2 _27677_ (.A(_07107_),
    .B(_07028_),
    .X(_11005_));
 sky130_fd_sc_hd__clkbuf_4 _27678_ (.A(_09152_),
    .X(_11006_));
 sky130_fd_sc_hd__nand3_4 _27679_ (.A(_11006_),
    .B(_07104_),
    .C(_06762_),
    .Y(_11007_));
 sky130_fd_sc_hd__buf_4 _27680_ (.A(_08627_),
    .X(_11008_));
 sky130_fd_sc_hd__clkbuf_4 _27681_ (.A(_09153_),
    .X(_11009_));
 sky130_fd_sc_hd__a22o_1 _27682_ (.A1(_11008_),
    .A2(_07481_),
    .B1(_11009_),
    .B2(_07034_),
    .X(_11010_));
 sky130_fd_sc_hd__o21ai_4 _27683_ (.A1(_08332_),
    .A2(_11007_),
    .B1(_11010_),
    .Y(_11011_));
 sky130_fd_sc_hd__xor2_4 _27684_ (.A(_11005_),
    .B(_11011_),
    .X(_11012_));
 sky130_fd_sc_hd__xnor2_4 _27685_ (.A(_11004_),
    .B(_11012_),
    .Y(_11013_));
 sky130_fd_sc_hd__xnor2_4 _27686_ (.A(_11003_),
    .B(_11013_),
    .Y(_11014_));
 sky130_fd_sc_hd__or2b_2 _27687_ (.A(_10868_),
    .B_N(_10863_),
    .X(_11015_));
 sky130_fd_sc_hd__o21ai_4 _27688_ (.A1(_10861_),
    .A2(_10869_),
    .B1(_11015_),
    .Y(_11016_));
 sky130_fd_sc_hd__and2_2 _27689_ (.A(_07359_),
    .B(_06578_),
    .X(_11017_));
 sky130_fd_sc_hd__buf_4 _27690_ (.A(_08396_),
    .X(_11018_));
 sky130_fd_sc_hd__nand3_4 _27691_ (.A(_11018_),
    .B(_13979_),
    .C(_06280_),
    .Y(_11019_));
 sky130_fd_sc_hd__clkbuf_4 _27692_ (.A(_08637_),
    .X(_11020_));
 sky130_fd_sc_hd__a22o_2 _27693_ (.A1(_13972_),
    .A2(_06438_),
    .B1(_11020_),
    .B2(_06432_),
    .X(_11021_));
 sky130_fd_sc_hd__o21ai_4 _27694_ (.A1(_14348_),
    .A2(_11019_),
    .B1(_11021_),
    .Y(_11022_));
 sky130_fd_sc_hd__xor2_4 _27695_ (.A(_11017_),
    .B(_11022_),
    .X(_11023_));
 sky130_fd_sc_hd__buf_6 _27696_ (.A(_13967_),
    .X(_11024_));
 sky130_fd_sc_hd__buf_6 _27697_ (.A(_09876_),
    .X(_11025_));
 sky130_fd_sc_hd__nand3b_4 _27698_ (.A_N(_10865_),
    .B(_11025_),
    .C(_08210_),
    .Y(_11026_));
 sky130_fd_sc_hd__o31ai_4 _27699_ (.A1(_11024_),
    .A2(_14368_),
    .A3(_10867_),
    .B1(_11026_),
    .Y(_11027_));
 sky130_fd_sc_hd__clkbuf_2 _27700_ (.A(_09172_),
    .X(_11028_));
 sky130_fd_sc_hd__and2_2 _27701_ (.A(_11028_),
    .B(_06285_),
    .X(_11029_));
 sky130_fd_sc_hd__clkbuf_4 _27702_ (.A(_13961_),
    .X(_11030_));
 sky130_fd_sc_hd__nand2_2 _27703_ (.A(_11030_),
    .B(_08720_),
    .Y(_11031_));
 sky130_fd_sc_hd__and2b_1 _27704_ (.A_N(_05699_),
    .B(_12805_),
    .X(_11032_));
 sky130_fd_sc_hd__xor2_4 _27705_ (.A(_11031_),
    .B(_11032_),
    .X(_11033_));
 sky130_fd_sc_hd__xor2_4 _27706_ (.A(_11029_),
    .B(_11033_),
    .X(_11034_));
 sky130_fd_sc_hd__xor2_4 _27707_ (.A(_11027_),
    .B(_11034_),
    .X(_11035_));
 sky130_fd_sc_hd__xor2_4 _27708_ (.A(_11023_),
    .B(_11035_),
    .X(_11036_));
 sky130_fd_sc_hd__xnor2_4 _27709_ (.A(_11016_),
    .B(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__xor2_4 _27710_ (.A(_11014_),
    .B(_11037_),
    .X(_11038_));
 sky130_fd_sc_hd__xnor2_1 _27711_ (.A(_11002_),
    .B(_11038_),
    .Y(_11039_));
 sky130_fd_sc_hd__or2b_2 _27712_ (.A(_11000_),
    .B_N(_11039_),
    .X(_11040_));
 sky130_fd_sc_hd__or2b_2 _27713_ (.A(_11039_),
    .B_N(_11000_),
    .X(_11041_));
 sky130_fd_sc_hd__a21o_1 _27714_ (.A1(_10872_),
    .A2(_10845_),
    .B1(_10874_),
    .X(_11042_));
 sky130_fd_sc_hd__a21o_1 _27715_ (.A1(_11040_),
    .A2(_11041_),
    .B1(_11042_),
    .X(_11043_));
 sky130_fd_sc_hd__nand3_4 _27716_ (.A(_11042_),
    .B(_11040_),
    .C(_11041_),
    .Y(_11044_));
 sky130_fd_sc_hd__and2b_1 _27717_ (.A_N(_10901_),
    .B(_10889_),
    .X(_11045_));
 sky130_fd_sc_hd__a21oi_4 _27718_ (.A1(_10900_),
    .A2(_10891_),
    .B1(_11045_),
    .Y(_11046_));
 sky130_fd_sc_hd__and2_1 _27719_ (.A(_10840_),
    .B(_10824_),
    .X(_11047_));
 sky130_fd_sc_hd__o21bai_2 _27720_ (.A1(_10822_),
    .A2(_10841_),
    .B1_N(_11047_),
    .Y(_11048_));
 sky130_fd_sc_hd__a2bb2oi_4 _27721_ (.A1_N(_14048_),
    .A2_N(_10885_),
    .B1(_10568_),
    .B2(_10884_),
    .Y(_11049_));
 sky130_fd_sc_hd__xor2_4 _27722_ (.A(_11049_),
    .B(_10414_),
    .X(_11050_));
 sky130_fd_sc_hd__inv_4 _27723_ (.A(_11050_),
    .Y(_11051_));
 sky130_fd_sc_hd__nor2_1 _27724_ (.A(_10893_),
    .B(_10898_),
    .Y(_11052_));
 sky130_fd_sc_hd__o21bai_4 _27725_ (.A1(_10892_),
    .A2(_10899_),
    .B1_N(_11052_),
    .Y(_11053_));
 sky130_fd_sc_hd__a2bb2oi_4 _27726_ (.A1_N(_14281_),
    .A2_N(_10895_),
    .B1(_10894_),
    .B2(_10896_),
    .Y(_11054_));
 sky130_fd_sc_hd__a2bb2oi_4 _27727_ (.A1_N(_14299_),
    .A2_N(_10828_),
    .B1(_10826_),
    .B2(_10830_),
    .Y(_11055_));
 sky130_fd_sc_hd__and2_1 _27728_ (.A(_12777_),
    .B(_06489_),
    .X(_11056_));
 sky130_fd_sc_hd__buf_6 _27729_ (.A(_11056_),
    .X(_11057_));
 sky130_fd_sc_hd__nand3_4 _27730_ (.A(_07295_),
    .B(_05815_),
    .C(_08806_),
    .Y(_11058_));
 sky130_fd_sc_hd__a22o_2 _27731_ (.A1(_07820_),
    .A2(_08165_),
    .B1(_05815_),
    .B2(_08171_),
    .X(_11059_));
 sky130_fd_sc_hd__o21ai_4 _27732_ (.A1(_14275_),
    .A2(_11058_),
    .B1(_11059_),
    .Y(_11060_));
 sky130_fd_sc_hd__xor2_4 _27733_ (.A(_11057_),
    .B(_11060_),
    .X(_11061_));
 sky130_fd_sc_hd__xnor2_4 _27734_ (.A(_11055_),
    .B(_11061_),
    .Y(_11062_));
 sky130_fd_sc_hd__xor2_4 _27735_ (.A(_11054_),
    .B(_11062_),
    .X(_11063_));
 sky130_fd_sc_hd__xnor2_4 _27736_ (.A(_11053_),
    .B(_11063_),
    .Y(_11064_));
 sky130_fd_sc_hd__xor2_4 _27737_ (.A(_11051_),
    .B(_11064_),
    .X(_11065_));
 sky130_fd_sc_hd__xnor2_2 _27738_ (.A(_11048_),
    .B(_11065_),
    .Y(_11066_));
 sky130_fd_sc_hd__xnor2_1 _27739_ (.A(_11046_),
    .B(_11066_),
    .Y(_11067_));
 sky130_fd_sc_hd__a21boi_1 _27740_ (.A1(_11043_),
    .A2(_11044_),
    .B1_N(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__nand3b_4 _27741_ (.A_N(_11067_),
    .B(_11043_),
    .C(_11044_),
    .Y(_11069_));
 sky130_vsdinv _27742_ (.A(_11069_),
    .Y(_11070_));
 sky130_fd_sc_hd__o21ai_4 _27743_ (.A1(_10904_),
    .A2(_10877_),
    .B1(_10879_),
    .Y(_11071_));
 sky130_fd_sc_hd__o21bai_1 _27744_ (.A1(_11068_),
    .A2(_11070_),
    .B1_N(_11071_),
    .Y(_11072_));
 sky130_fd_sc_hd__a21bo_2 _27745_ (.A1(_11043_),
    .A2(_11044_),
    .B1_N(_11067_),
    .X(_11073_));
 sky130_fd_sc_hd__nand3_4 _27746_ (.A(_11073_),
    .B(_11069_),
    .C(_11071_),
    .Y(_11074_));
 sky130_fd_sc_hd__nand2_2 _27747_ (.A(_10902_),
    .B(_10883_),
    .Y(_11075_));
 sky130_fd_sc_hd__or2_2 _27748_ (.A(_10881_),
    .B(_10903_),
    .X(_11076_));
 sky130_fd_sc_hd__nand3b_2 _27749_ (.A_N(_10731_),
    .B(_14038_),
    .C(_05442_),
    .Y(_11077_));
 sky130_fd_sc_hd__a21boi_4 _27750_ (.A1(_10888_),
    .A2(_10414_),
    .B1_N(_11077_),
    .Y(_11078_));
 sky130_fd_sc_hd__nand3_4 _27751_ (.A(_10609_),
    .B(_10135_),
    .C(_10610_),
    .Y(_11079_));
 sky130_fd_sc_hd__o21ai_2 _27752_ (.A1(_10609_),
    .A2(_10764_),
    .B1(_11079_),
    .Y(_11080_));
 sky130_fd_sc_hd__xnor2_2 _27753_ (.A(_11078_),
    .B(_11080_),
    .Y(_11081_));
 sky130_fd_sc_hd__and2_1 _27754_ (.A(_10916_),
    .B(_10913_),
    .X(_11082_));
 sky130_fd_sc_hd__a21o_1 _27755_ (.A1(_10612_),
    .A2(_10915_),
    .B1(_11082_),
    .X(_11083_));
 sky130_fd_sc_hd__xor2_2 _27756_ (.A(_11081_),
    .B(_11083_),
    .X(_11084_));
 sky130_fd_sc_hd__xor2_1 _27757_ (.A(_09985_),
    .B(_11084_),
    .X(_11085_));
 sky130_fd_sc_hd__a21bo_2 _27758_ (.A1(_11075_),
    .A2(_11076_),
    .B1_N(_11085_),
    .X(_11086_));
 sky130_fd_sc_hd__nand3b_4 _27759_ (.A_N(_11085_),
    .B(_11075_),
    .C(_11076_),
    .Y(_11087_));
 sky130_fd_sc_hd__o21ba_1 _27760_ (.A1(_10446_),
    .A2(_10920_),
    .B1_N(_10921_),
    .X(_11088_));
 sky130_vsdinv _27761_ (.A(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__a21o_1 _27762_ (.A1(_11086_),
    .A2(_11087_),
    .B1(_11089_),
    .X(_11090_));
 sky130_fd_sc_hd__nand3_4 _27763_ (.A(_11086_),
    .B(_11089_),
    .C(_11087_),
    .Y(_11091_));
 sky130_fd_sc_hd__nand2_4 _27764_ (.A(_11090_),
    .B(_11091_),
    .Y(_11092_));
 sky130_fd_sc_hd__a21boi_1 _27765_ (.A1(_11072_),
    .A2(_11074_),
    .B1_N(_11092_),
    .Y(_11093_));
 sky130_fd_sc_hd__a21oi_4 _27766_ (.A1(_11073_),
    .A2(_11069_),
    .B1(_11071_),
    .Y(_11094_));
 sky130_vsdinv _27767_ (.A(_11074_),
    .Y(_11095_));
 sky130_fd_sc_hd__nor3_4 _27768_ (.A(_11092_),
    .B(_11094_),
    .C(_11095_),
    .Y(_11096_));
 sky130_fd_sc_hd__o21ai_2 _27769_ (.A1(_10935_),
    .A2(_10936_),
    .B1(_10912_),
    .Y(_11097_));
 sky130_fd_sc_hd__o21bai_2 _27770_ (.A1(_11093_),
    .A2(_11096_),
    .B1_N(_11097_),
    .Y(_11098_));
 sky130_fd_sc_hd__o21ai_2 _27771_ (.A1(_11094_),
    .A2(_11095_),
    .B1(_11092_),
    .Y(_11099_));
 sky130_fd_sc_hd__nand3b_2 _27772_ (.A_N(_11092_),
    .B(_11074_),
    .C(_11072_),
    .Y(_11100_));
 sky130_fd_sc_hd__nand3_4 _27773_ (.A(_11099_),
    .B(_11100_),
    .C(_11097_),
    .Y(_11101_));
 sky130_fd_sc_hd__a21boi_4 _27774_ (.A1(_10930_),
    .A2(_10927_),
    .B1_N(_10926_),
    .Y(_11102_));
 sky130_fd_sc_hd__xor2_4 _27775_ (.A(_10325_),
    .B(_11102_),
    .X(_11103_));
 sky130_fd_sc_hd__a21oi_1 _27776_ (.A1(_11098_),
    .A2(_11101_),
    .B1(_11103_),
    .Y(_11104_));
 sky130_fd_sc_hd__nand3_4 _27777_ (.A(_11098_),
    .B(_11103_),
    .C(_11101_),
    .Y(_11105_));
 sky130_vsdinv _27778_ (.A(_11105_),
    .Y(_11106_));
 sky130_fd_sc_hd__o21ai_4 _27779_ (.A1(_10948_),
    .A2(_10949_),
    .B1(_10944_),
    .Y(_11107_));
 sky130_fd_sc_hd__o21bai_2 _27780_ (.A1(_11104_),
    .A2(_11106_),
    .B1_N(_11107_),
    .Y(_11108_));
 sky130_fd_sc_hd__nand2_1 _27781_ (.A(_11098_),
    .B(_11101_),
    .Y(_11109_));
 sky130_vsdinv _27782_ (.A(_11103_),
    .Y(_11110_));
 sky130_fd_sc_hd__nand2_2 _27783_ (.A(_11109_),
    .B(_11110_),
    .Y(_11111_));
 sky130_fd_sc_hd__nand3_4 _27784_ (.A(_11111_),
    .B(_11105_),
    .C(_11107_),
    .Y(_11112_));
 sky130_fd_sc_hd__and2_2 _27785_ (.A(_10945_),
    .B(_10178_),
    .X(_11113_));
 sky130_fd_sc_hd__a21oi_1 _27786_ (.A1(_11108_),
    .A2(_11112_),
    .B1(_11113_),
    .Y(_11114_));
 sky130_vsdinv _27787_ (.A(_11113_),
    .Y(_11115_));
 sky130_fd_sc_hd__a21oi_2 _27788_ (.A1(_11111_),
    .A2(_11105_),
    .B1(_11107_),
    .Y(_11116_));
 sky130_fd_sc_hd__nor3b_4 _27789_ (.A(_11115_),
    .B(_11116_),
    .C_N(_11112_),
    .Y(_11117_));
 sky130_fd_sc_hd__o21ai_2 _27790_ (.A1(_10961_),
    .A2(_10962_),
    .B1(_10959_),
    .Y(_11118_));
 sky130_fd_sc_hd__o21bai_2 _27791_ (.A1(_11114_),
    .A2(_11117_),
    .B1_N(_11118_),
    .Y(_11119_));
 sky130_fd_sc_hd__a21o_1 _27792_ (.A1(_11108_),
    .A2(_11112_),
    .B1(_11113_),
    .X(_11120_));
 sky130_fd_sc_hd__nand3_2 _27793_ (.A(_11108_),
    .B(_11113_),
    .C(_11112_),
    .Y(_11121_));
 sky130_fd_sc_hd__nand3_4 _27794_ (.A(_11120_),
    .B(_11118_),
    .C(_11121_),
    .Y(_11122_));
 sky130_fd_sc_hd__and2_1 _27795_ (.A(_11119_),
    .B(_11122_),
    .X(_11123_));
 sky130_fd_sc_hd__o21ai_1 _27796_ (.A1(_10973_),
    .A2(_10978_),
    .B1(_10972_),
    .Y(_11124_));
 sky130_fd_sc_hd__xor2_1 _27797_ (.A(_11123_),
    .B(_11124_),
    .X(_02666_));
 sky130_fd_sc_hd__nor2_1 _27798_ (.A(_10989_),
    .B(_10996_),
    .Y(_11125_));
 sky130_fd_sc_hd__o21ba_1 _27799_ (.A1(_10988_),
    .A2(_10997_),
    .B1_N(_11125_),
    .X(_11126_));
 sky130_fd_sc_hd__nor2_1 _27800_ (.A(_11004_),
    .B(_11012_),
    .Y(_11127_));
 sky130_fd_sc_hd__o21bai_1 _27801_ (.A1(_11003_),
    .A2(_11013_),
    .B1_N(_11127_),
    .Y(_11128_));
 sky130_fd_sc_hd__a2bb2oi_4 _27802_ (.A1_N(_14311_),
    .A2_N(_10993_),
    .B1(_10990_),
    .B2(_10994_),
    .Y(_11129_));
 sky130_fd_sc_hd__and2_2 _27803_ (.A(_06472_),
    .B(_10829_),
    .X(_11130_));
 sky130_fd_sc_hd__nand3_4 _27804_ (.A(_10991_),
    .B(_10992_),
    .C(_07575_),
    .Y(_11131_));
 sky130_fd_sc_hd__buf_4 _27805_ (.A(_09197_),
    .X(_11132_));
 sky130_fd_sc_hd__buf_4 _27806_ (.A(_08864_),
    .X(_11133_));
 sky130_fd_sc_hd__a22o_2 _27807_ (.A1(_11132_),
    .A2(_08885_),
    .B1(_11133_),
    .B2(_07775_),
    .X(_11134_));
 sky130_fd_sc_hd__o21ai_4 _27808_ (.A1(_14304_),
    .A2(_11131_),
    .B1(_11134_),
    .Y(_11135_));
 sky130_fd_sc_hd__xor2_4 _27809_ (.A(_11130_),
    .B(_11135_),
    .X(_11136_));
 sky130_fd_sc_hd__xnor2_2 _27810_ (.A(_11129_),
    .B(_11136_),
    .Y(_11137_));
 sky130_fd_sc_hd__buf_2 _27811_ (.A(_08806_),
    .X(_11138_));
 sky130_fd_sc_hd__and2_2 _27812_ (.A(_06061_),
    .B(_11138_),
    .X(_11139_));
 sky130_fd_sc_hd__or4_4 _27813_ (.A(_14011_),
    .B(_14016_),
    .C(_14286_),
    .D(_14292_),
    .X(_11140_));
 sky130_fd_sc_hd__a22o_1 _27814_ (.A1(_10984_),
    .A2(_10825_),
    .B1(_10705_),
    .B2(_08489_),
    .X(_11141_));
 sky130_fd_sc_hd__nand2_2 _27815_ (.A(_11140_),
    .B(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__xor2_4 _27816_ (.A(_11139_),
    .B(_11142_),
    .X(_11143_));
 sky130_fd_sc_hd__xor2_2 _27817_ (.A(_11137_),
    .B(_11143_),
    .X(_11144_));
 sky130_fd_sc_hd__xnor2_1 _27818_ (.A(_11128_),
    .B(_11144_),
    .Y(_11145_));
 sky130_fd_sc_hd__xor2_1 _27819_ (.A(_11126_),
    .B(_11145_),
    .X(_11146_));
 sky130_vsdinv _27820_ (.A(_11146_),
    .Y(_11147_));
 sky130_fd_sc_hd__and2_1 _27821_ (.A(_11036_),
    .B(_11016_),
    .X(_11148_));
 sky130_fd_sc_hd__o21bai_4 _27822_ (.A1(_11014_),
    .A2(_11037_),
    .B1_N(_11148_),
    .Y(_11149_));
 sky130_fd_sc_hd__a2bb2oi_1 _27823_ (.A1_N(_14329_),
    .A2_N(_11007_),
    .B1(_11005_),
    .B2(_11010_),
    .Y(_11150_));
 sky130_vsdinv _27824_ (.A(_11150_),
    .Y(_11151_));
 sky130_fd_sc_hd__a2bb2oi_4 _27825_ (.A1_N(_14348_),
    .A2_N(_11019_),
    .B1(_11017_),
    .B2(_11021_),
    .Y(_11152_));
 sky130_fd_sc_hd__and2_4 _27826_ (.A(_08400_),
    .B(_08085_),
    .X(_11153_));
 sky130_fd_sc_hd__nand3_4 _27827_ (.A(_09152_),
    .B(_09153_),
    .C(_08701_),
    .Y(_11154_));
 sky130_fd_sc_hd__a22o_2 _27828_ (.A1(_08627_),
    .A2(_06940_),
    .B1(_08628_),
    .B2(_07036_),
    .X(_11155_));
 sky130_fd_sc_hd__o21ai_4 _27829_ (.A1(_08699_),
    .A2(_11154_),
    .B1(_11155_),
    .Y(_11156_));
 sky130_fd_sc_hd__xor2_4 _27830_ (.A(_11153_),
    .B(_11156_),
    .X(_11157_));
 sky130_fd_sc_hd__xnor2_4 _27831_ (.A(_11152_),
    .B(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__xor2_4 _27832_ (.A(_11151_),
    .B(_11158_),
    .X(_11159_));
 sky130_fd_sc_hd__or2b_1 _27833_ (.A(_11034_),
    .B_N(_11027_),
    .X(_11160_));
 sky130_fd_sc_hd__o21ai_4 _27834_ (.A1(_11023_),
    .A2(_11035_),
    .B1(_11160_),
    .Y(_11161_));
 sky130_fd_sc_hd__clkbuf_2 _27835_ (.A(_07873_),
    .X(_11162_));
 sky130_fd_sc_hd__and2_2 _27836_ (.A(_11162_),
    .B(_06762_),
    .X(_11163_));
 sky130_fd_sc_hd__buf_6 _27837_ (.A(_11020_),
    .X(_11164_));
 sky130_fd_sc_hd__nand3_4 _27838_ (.A(_13973_),
    .B(_11164_),
    .C(_06432_),
    .Y(_11165_));
 sky130_fd_sc_hd__buf_4 _27839_ (.A(_13978_),
    .X(_11166_));
 sky130_fd_sc_hd__a22o_2 _27840_ (.A1(_11018_),
    .A2(_06432_),
    .B1(_11166_),
    .B2(_06578_),
    .X(_11167_));
 sky130_fd_sc_hd__o21ai_4 _27841_ (.A1(_14342_),
    .A2(_11165_),
    .B1(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__xor2_4 _27842_ (.A(_11163_),
    .B(_11168_),
    .X(_11169_));
 sky130_fd_sc_hd__nand3b_4 _27843_ (.A_N(_11031_),
    .B(_11025_),
    .C(_14374_),
    .Y(_11170_));
 sky130_fd_sc_hd__o31ai_4 _27844_ (.A1(_13968_),
    .A2(_14361_),
    .A3(_11033_),
    .B1(_11170_),
    .Y(_11171_));
 sky130_fd_sc_hd__and2_2 _27845_ (.A(_07946_),
    .B(_06438_),
    .X(_11172_));
 sky130_fd_sc_hd__nand2_2 _27846_ (.A(_11030_),
    .B(_05913_),
    .Y(_11173_));
 sky130_fd_sc_hd__and2b_1 _27847_ (.A_N(_08720_),
    .B(_09025_),
    .X(_11174_));
 sky130_fd_sc_hd__xor2_4 _27848_ (.A(_11173_),
    .B(_11174_),
    .X(_11175_));
 sky130_fd_sc_hd__xor2_4 _27849_ (.A(_11172_),
    .B(_11175_),
    .X(_11176_));
 sky130_fd_sc_hd__xor2_4 _27850_ (.A(_11171_),
    .B(_11176_),
    .X(_11177_));
 sky130_fd_sc_hd__xor2_4 _27851_ (.A(_11169_),
    .B(_11177_),
    .X(_11178_));
 sky130_fd_sc_hd__xnor2_4 _27852_ (.A(_11161_),
    .B(_11178_),
    .Y(_11179_));
 sky130_fd_sc_hd__xor2_4 _27853_ (.A(_11159_),
    .B(_11179_),
    .X(_11180_));
 sky130_fd_sc_hd__xnor2_4 _27854_ (.A(_11149_),
    .B(_11180_),
    .Y(_11181_));
 sky130_fd_sc_hd__xor2_4 _27855_ (.A(_11147_),
    .B(_11181_),
    .X(_11182_));
 sky130_fd_sc_hd__a21bo_1 _27856_ (.A1(_11038_),
    .A2(_11002_),
    .B1_N(_11041_),
    .X(_11183_));
 sky130_fd_sc_hd__nor2_2 _27857_ (.A(_11182_),
    .B(_11183_),
    .Y(_11184_));
 sky130_vsdinv _27858_ (.A(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__nand2_2 _27859_ (.A(_11183_),
    .B(_11182_),
    .Y(_11186_));
 sky130_fd_sc_hd__clkbuf_4 _27860_ (.A(_11051_),
    .X(_11187_));
 sky130_fd_sc_hd__nand2_1 _27861_ (.A(_11063_),
    .B(_11053_),
    .Y(_11188_));
 sky130_fd_sc_hd__o21a_2 _27862_ (.A1(_11187_),
    .A2(_11064_),
    .B1(_11188_),
    .X(_11189_));
 sky130_fd_sc_hd__and2_1 _27863_ (.A(_10998_),
    .B(_10982_),
    .X(_11190_));
 sky130_fd_sc_hd__o21bai_4 _27864_ (.A1(_10980_),
    .A2(_10999_),
    .B1_N(_11190_),
    .Y(_11191_));
 sky130_fd_sc_hd__nor2_1 _27865_ (.A(_11055_),
    .B(_11061_),
    .Y(_11192_));
 sky130_fd_sc_hd__o21bai_4 _27866_ (.A1(_11054_),
    .A2(_11062_),
    .B1_N(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__a2bb2oi_4 _27867_ (.A1_N(_14277_),
    .A2_N(_11058_),
    .B1(_11057_),
    .B2(_11059_),
    .Y(_11194_));
 sky130_fd_sc_hd__a2bb2oi_4 _27868_ (.A1_N(_14293_),
    .A2_N(_10985_),
    .B1(_10983_),
    .B2(_10986_),
    .Y(_11195_));
 sky130_fd_sc_hd__nand2_4 _27869_ (.A(_07820_),
    .B(_08595_),
    .Y(_11196_));
 sky130_fd_sc_hd__nand2_4 _27870_ (.A(_09283_),
    .B(_05815_),
    .Y(_11197_));
 sky130_fd_sc_hd__xnor2_4 _27871_ (.A(_11196_),
    .B(_11197_),
    .Y(_11198_));
 sky130_fd_sc_hd__xor2_4 _27872_ (.A(_11057_),
    .B(_11198_),
    .X(_11199_));
 sky130_fd_sc_hd__xnor2_4 _27873_ (.A(_11195_),
    .B(_11199_),
    .Y(_11200_));
 sky130_fd_sc_hd__xor2_4 _27874_ (.A(_11194_),
    .B(_11200_),
    .X(_11201_));
 sky130_fd_sc_hd__xnor2_4 _27875_ (.A(_11193_),
    .B(_11201_),
    .Y(_11202_));
 sky130_fd_sc_hd__xor2_4 _27876_ (.A(_11051_),
    .B(_11202_),
    .X(_11203_));
 sky130_fd_sc_hd__xnor2_4 _27877_ (.A(_11191_),
    .B(_11203_),
    .Y(_11204_));
 sky130_fd_sc_hd__xor2_4 _27878_ (.A(_11189_),
    .B(_11204_),
    .X(_11205_));
 sky130_fd_sc_hd__a21oi_1 _27879_ (.A1(_11185_),
    .A2(_11186_),
    .B1(_11205_),
    .Y(_11206_));
 sky130_fd_sc_hd__nand3b_4 _27880_ (.A_N(_11184_),
    .B(_11205_),
    .C(_11186_),
    .Y(_11207_));
 sky130_vsdinv _27881_ (.A(_11207_),
    .Y(_11208_));
 sky130_fd_sc_hd__nand2_2 _27882_ (.A(_11069_),
    .B(_11044_),
    .Y(_11209_));
 sky130_fd_sc_hd__o21bai_2 _27883_ (.A1(_11206_),
    .A2(_11208_),
    .B1_N(_11209_),
    .Y(_11210_));
 sky130_fd_sc_hd__a21o_1 _27884_ (.A1(_11185_),
    .A2(_11186_),
    .B1(_11205_),
    .X(_11211_));
 sky130_fd_sc_hd__nand3_4 _27885_ (.A(_11211_),
    .B(_11207_),
    .C(_11209_),
    .Y(_11212_));
 sky130_fd_sc_hd__or2b_1 _27886_ (.A(_11081_),
    .B_N(_11083_),
    .X(_11213_));
 sky130_fd_sc_hd__o21a_2 _27887_ (.A1(_10446_),
    .A2(_11084_),
    .B1(_11213_),
    .X(_11214_));
 sky130_fd_sc_hd__a21boi_4 _27888_ (.A1(_10414_),
    .A2(_11049_),
    .B1_N(_11077_),
    .Y(_11215_));
 sky130_fd_sc_hd__o31ai_1 _27889_ (.A1(_10135_),
    .A2(_10609_),
    .A3(_10610_),
    .B1(_11078_),
    .Y(_11216_));
 sky130_fd_sc_hd__and2_1 _27890_ (.A(_11216_),
    .B(_11079_),
    .X(_11217_));
 sky130_fd_sc_hd__xor2_4 _27891_ (.A(_11215_),
    .B(_11217_),
    .X(_11218_));
 sky130_fd_sc_hd__xor2_4 _27892_ (.A(_11218_),
    .B(_09978_),
    .X(_11219_));
 sky130_fd_sc_hd__nand2_1 _27893_ (.A(_11065_),
    .B(_11048_),
    .Y(_11220_));
 sky130_fd_sc_hd__o21ai_4 _27894_ (.A1(_11046_),
    .A2(_11066_),
    .B1(_11220_),
    .Y(_11221_));
 sky130_fd_sc_hd__xnor2_4 _27895_ (.A(_11219_),
    .B(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__xnor2_2 _27896_ (.A(_11214_),
    .B(_11222_),
    .Y(_11223_));
 sky130_fd_sc_hd__a21bo_1 _27897_ (.A1(_11210_),
    .A2(_11212_),
    .B1_N(_11223_),
    .X(_11224_));
 sky130_fd_sc_hd__nand3b_4 _27898_ (.A_N(_11223_),
    .B(_11210_),
    .C(_11212_),
    .Y(_11225_));
 sky130_fd_sc_hd__o21ai_4 _27899_ (.A1(_11092_),
    .A2(_11094_),
    .B1(_11074_),
    .Y(_11226_));
 sky130_fd_sc_hd__a21oi_2 _27900_ (.A1(_11224_),
    .A2(_11225_),
    .B1(_11226_),
    .Y(_11227_));
 sky130_fd_sc_hd__nand3_4 _27901_ (.A(_11224_),
    .B(_11225_),
    .C(_11226_),
    .Y(_11228_));
 sky130_vsdinv _27902_ (.A(_11228_),
    .Y(_11229_));
 sky130_fd_sc_hd__a21boi_4 _27903_ (.A1(_11089_),
    .A2(_11087_),
    .B1_N(_11086_),
    .Y(_11230_));
 sky130_fd_sc_hd__xor2_4 _27904_ (.A(net413),
    .B(_11230_),
    .X(_11231_));
 sky130_fd_sc_hd__o21bai_2 _27905_ (.A1(_11227_),
    .A2(_11229_),
    .B1_N(_11231_),
    .Y(_11232_));
 sky130_fd_sc_hd__a21boi_1 _27906_ (.A1(_11210_),
    .A2(_11212_),
    .B1_N(_11223_),
    .Y(_11233_));
 sky130_vsdinv _27907_ (.A(_11225_),
    .Y(_11234_));
 sky130_fd_sc_hd__o21bai_2 _27908_ (.A1(_11233_),
    .A2(_11234_),
    .B1_N(_11226_),
    .Y(_11235_));
 sky130_fd_sc_hd__nand3_4 _27909_ (.A(_11235_),
    .B(_11231_),
    .C(_11228_),
    .Y(_11236_));
 sky130_fd_sc_hd__nand2_2 _27910_ (.A(_11105_),
    .B(_11101_),
    .Y(_11237_));
 sky130_fd_sc_hd__nand3_4 _27911_ (.A(_11232_),
    .B(_11236_),
    .C(_11237_),
    .Y(_11238_));
 sky130_fd_sc_hd__a21oi_1 _27912_ (.A1(_11235_),
    .A2(_11228_),
    .B1(_11231_),
    .Y(_11239_));
 sky130_vsdinv _27913_ (.A(_11236_),
    .Y(_11240_));
 sky130_fd_sc_hd__o21bai_2 _27914_ (.A1(_11239_),
    .A2(_11240_),
    .B1_N(_11237_),
    .Y(_11241_));
 sky130_fd_sc_hd__buf_4 _27915_ (.A(_10812_),
    .X(_11242_));
 sky130_fd_sc_hd__buf_4 _27916_ (.A(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__o2bb2ai_2 _27917_ (.A1_N(_11238_),
    .A2_N(_11241_),
    .B1(_11243_),
    .B2(_11102_),
    .Y(_11244_));
 sky130_fd_sc_hd__a21oi_4 _27918_ (.A1(_10932_),
    .A2(_10926_),
    .B1(_10813_),
    .Y(_11245_));
 sky130_fd_sc_hd__nand3_4 _27919_ (.A(_11241_),
    .B(_11245_),
    .C(_11238_),
    .Y(_11246_));
 sky130_fd_sc_hd__a21boi_1 _27920_ (.A1(_11108_),
    .A2(_11113_),
    .B1_N(_11112_),
    .Y(_11247_));
 sky130_vsdinv _27921_ (.A(_11247_),
    .Y(_11248_));
 sky130_fd_sc_hd__a21o_1 _27922_ (.A1(_11244_),
    .A2(_11246_),
    .B1(_11248_),
    .X(_11249_));
 sky130_fd_sc_hd__nand3_4 _27923_ (.A(_11244_),
    .B(_11246_),
    .C(_11248_),
    .Y(_11250_));
 sky130_fd_sc_hd__nand2_2 _27924_ (.A(_11249_),
    .B(_11250_),
    .Y(_11251_));
 sky130_fd_sc_hd__nand2_1 _27925_ (.A(_11119_),
    .B(_11122_),
    .Y(_11252_));
 sky130_fd_sc_hd__nor2_1 _27926_ (.A(_10973_),
    .B(_11252_),
    .Y(_11253_));
 sky130_fd_sc_hd__nand2_1 _27927_ (.A(_10975_),
    .B(_11253_),
    .Y(_11254_));
 sky130_fd_sc_hd__nor2_1 _27928_ (.A(_10661_),
    .B(_11254_),
    .Y(_11255_));
 sky130_fd_sc_hd__nand3_2 _27929_ (.A(_08567_),
    .B(_10030_),
    .C(_11255_),
    .Y(_11256_));
 sky130_fd_sc_hd__nand2_1 _27930_ (.A(_10036_),
    .B(_11255_),
    .Y(_11257_));
 sky130_fd_sc_hd__a21oi_1 _27931_ (.A1(_10647_),
    .A2(_10643_),
    .B1(_10642_),
    .Y(_11258_));
 sky130_fd_sc_hd__nor3_2 _27932_ (.A(_11258_),
    .B(_10806_),
    .C(_10808_),
    .Y(_11259_));
 sky130_fd_sc_hd__nor2_1 _27933_ (.A(_10976_),
    .B(_11259_),
    .Y(_11260_));
 sky130_fd_sc_hd__nand2_1 _27934_ (.A(_10654_),
    .B(_11260_),
    .Y(_11261_));
 sky130_fd_sc_hd__and2_1 _27935_ (.A(_10969_),
    .B(_10972_),
    .X(_11262_));
 sky130_fd_sc_hd__nand2_1 _27936_ (.A(_11123_),
    .B(_11262_),
    .Y(_11263_));
 sky130_fd_sc_hd__nor2_2 _27937_ (.A(_11261_),
    .B(_11263_),
    .Y(_11264_));
 sky130_fd_sc_hd__nand3_2 _27938_ (.A(_11123_),
    .B(_11262_),
    .C(_10977_),
    .Y(_11265_));
 sky130_fd_sc_hd__or2b_1 _27939_ (.A(_10972_),
    .B_N(_11119_),
    .X(_11266_));
 sky130_fd_sc_hd__nand3_4 _27940_ (.A(_11265_),
    .B(_11122_),
    .C(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__a21oi_4 _27941_ (.A1(_11264_),
    .A2(_10665_),
    .B1(_11267_),
    .Y(_11268_));
 sky130_fd_sc_hd__nand3_4 _27942_ (.A(_11256_),
    .B(_11257_),
    .C(_11268_),
    .Y(_11269_));
 sky130_fd_sc_hd__xnor2_1 _27943_ (.A(_11251_),
    .B(_11269_),
    .Y(_02667_));
 sky130_fd_sc_hd__and2_1 _27944_ (.A(_11180_),
    .B(_11149_),
    .X(_11270_));
 sky130_fd_sc_hd__o21ba_1 _27945_ (.A1(_11147_),
    .A2(_11181_),
    .B1_N(_11270_),
    .X(_11271_));
 sky130_fd_sc_hd__nor2_1 _27946_ (.A(_11129_),
    .B(_11136_),
    .Y(_11272_));
 sky130_fd_sc_hd__o21ba_1 _27947_ (.A1(_11137_),
    .A2(_11143_),
    .B1_N(_11272_),
    .X(_11273_));
 sky130_fd_sc_hd__or2b_1 _27948_ (.A(_11158_),
    .B_N(_11151_),
    .X(_11274_));
 sky130_fd_sc_hd__o21ai_2 _27949_ (.A1(_11152_),
    .A2(_11157_),
    .B1(_11274_),
    .Y(_11275_));
 sky130_fd_sc_hd__a2bb2oi_4 _27950_ (.A1_N(_14305_),
    .A2_N(_11131_),
    .B1(_11130_),
    .B2(_11134_),
    .Y(_11276_));
 sky130_fd_sc_hd__and2_2 _27951_ (.A(_09388_),
    .B(_08064_),
    .X(_11277_));
 sky130_fd_sc_hd__nand3_4 _27952_ (.A(_11132_),
    .B(_11133_),
    .C(_07569_),
    .Y(_11278_));
 sky130_fd_sc_hd__a22o_2 _27953_ (.A1(_10515_),
    .A2(_07477_),
    .B1(_10516_),
    .B2(_07578_),
    .X(_11279_));
 sky130_fd_sc_hd__o21ai_4 _27954_ (.A1(_14298_),
    .A2(_11278_),
    .B1(_11279_),
    .Y(_11280_));
 sky130_fd_sc_hd__xor2_4 _27955_ (.A(_11277_),
    .B(_11280_),
    .X(_11281_));
 sky130_fd_sc_hd__xnor2_2 _27956_ (.A(_11276_),
    .B(_11281_),
    .Y(_11282_));
 sky130_fd_sc_hd__and2_2 _27957_ (.A(_06061_),
    .B(_08596_),
    .X(_11283_));
 sky130_fd_sc_hd__or4_4 _27958_ (.A(_14011_),
    .B(_14016_),
    .C(_14280_),
    .D(_14286_),
    .X(_11284_));
 sky130_fd_sc_hd__a22o_1 _27959_ (.A1(_10984_),
    .A2(_08157_),
    .B1(_10705_),
    .B2(_11138_),
    .X(_11285_));
 sky130_fd_sc_hd__nand2_2 _27960_ (.A(_11284_),
    .B(_11285_),
    .Y(_11286_));
 sky130_fd_sc_hd__xor2_4 _27961_ (.A(_11283_),
    .B(_11286_),
    .X(_11287_));
 sky130_fd_sc_hd__xor2_2 _27962_ (.A(_11282_),
    .B(_11287_),
    .X(_11288_));
 sky130_fd_sc_hd__xnor2_1 _27963_ (.A(_11275_),
    .B(_11288_),
    .Y(_11289_));
 sky130_fd_sc_hd__xor2_1 _27964_ (.A(_11273_),
    .B(_11289_),
    .X(_11290_));
 sky130_vsdinv _27965_ (.A(_11290_),
    .Y(_11291_));
 sky130_fd_sc_hd__and2_1 _27966_ (.A(_11178_),
    .B(_11161_),
    .X(_11292_));
 sky130_fd_sc_hd__o21bai_2 _27967_ (.A1(_11159_),
    .A2(_11179_),
    .B1_N(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__a2bb2oi_4 _27968_ (.A1_N(_14322_),
    .A2_N(_11154_),
    .B1(_11153_),
    .B2(_11155_),
    .Y(_11294_));
 sky130_fd_sc_hd__a2bb2oi_4 _27969_ (.A1_N(_14342_),
    .A2_N(_11165_),
    .B1(_11163_),
    .B2(_11167_),
    .Y(_11295_));
 sky130_fd_sc_hd__and2_2 _27970_ (.A(_07107_),
    .B(_07468_),
    .X(_11296_));
 sky130_fd_sc_hd__nand3_4 _27971_ (.A(_11008_),
    .B(_07104_),
    .C(_07028_),
    .Y(_11297_));
 sky130_fd_sc_hd__a22o_2 _27972_ (.A1(_11008_),
    .A2(_08330_),
    .B1(_11009_),
    .B2(_07473_),
    .X(_11298_));
 sky130_fd_sc_hd__o21ai_4 _27973_ (.A1(_08464_),
    .A2(_11297_),
    .B1(_11298_),
    .Y(_11299_));
 sky130_fd_sc_hd__xor2_4 _27974_ (.A(_11296_),
    .B(_11299_),
    .X(_11300_));
 sky130_fd_sc_hd__xnor2_4 _27975_ (.A(_11295_),
    .B(_11300_),
    .Y(_11301_));
 sky130_fd_sc_hd__xnor2_4 _27976_ (.A(_11294_),
    .B(_11301_),
    .Y(_11302_));
 sky130_fd_sc_hd__or2b_2 _27977_ (.A(_11176_),
    .B_N(_11171_),
    .X(_11303_));
 sky130_fd_sc_hd__o21ai_4 _27978_ (.A1(_11169_),
    .A2(_11177_),
    .B1(_11303_),
    .Y(_11304_));
 sky130_fd_sc_hd__and2_2 _27979_ (.A(_11162_),
    .B(_06941_),
    .X(_11305_));
 sky130_fd_sc_hd__nand3_4 _27980_ (.A(_11018_),
    .B(_11166_),
    .C(_06578_),
    .Y(_11306_));
 sky130_fd_sc_hd__a22o_2 _27981_ (.A1(_08397_),
    .A2(_06578_),
    .B1(_11020_),
    .B2(_07481_),
    .X(_11307_));
 sky130_fd_sc_hd__o21ai_4 _27982_ (.A1(_14334_),
    .A2(_11306_),
    .B1(_11307_),
    .Y(_11308_));
 sky130_fd_sc_hd__xor2_4 _27983_ (.A(_11305_),
    .B(_11308_),
    .X(_11309_));
 sky130_fd_sc_hd__nand3b_4 _27984_ (.A_N(_11173_),
    .B(_11025_),
    .C(_14367_),
    .Y(_11310_));
 sky130_fd_sc_hd__o31ai_4 _27985_ (.A1(_11024_),
    .A2(_14354_),
    .A3(_11175_),
    .B1(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__and2_2 _27986_ (.A(_11028_),
    .B(_06584_),
    .X(_11312_));
 sky130_fd_sc_hd__nand2_2 _27987_ (.A(_11030_),
    .B(_06155_),
    .Y(_11313_));
 sky130_fd_sc_hd__and2b_1 _27988_ (.A_N(_07650_),
    .B(_12805_),
    .X(_11314_));
 sky130_fd_sc_hd__xor2_4 _27989_ (.A(_11313_),
    .B(_11314_),
    .X(_11315_));
 sky130_fd_sc_hd__xor2_4 _27990_ (.A(_11312_),
    .B(_11315_),
    .X(_11316_));
 sky130_fd_sc_hd__xor2_4 _27991_ (.A(_11311_),
    .B(_11316_),
    .X(_11317_));
 sky130_fd_sc_hd__xor2_4 _27992_ (.A(_11309_),
    .B(_11317_),
    .X(_11318_));
 sky130_fd_sc_hd__xnor2_4 _27993_ (.A(_11304_),
    .B(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__xor2_4 _27994_ (.A(_11302_),
    .B(_11319_),
    .X(_11320_));
 sky130_fd_sc_hd__xnor2_2 _27995_ (.A(_11293_),
    .B(_11320_),
    .Y(_11321_));
 sky130_fd_sc_hd__xor2_2 _27996_ (.A(_11291_),
    .B(_11321_),
    .X(_11322_));
 sky130_fd_sc_hd__and2b_1 _27997_ (.A_N(_11271_),
    .B(_11322_),
    .X(_11323_));
 sky130_vsdinv _27998_ (.A(_11323_),
    .Y(_11324_));
 sky130_fd_sc_hd__or2b_2 _27999_ (.A(_11322_),
    .B_N(_11271_),
    .X(_11325_));
 sky130_fd_sc_hd__nand2_1 _28000_ (.A(_11201_),
    .B(_11193_),
    .Y(_11326_));
 sky130_fd_sc_hd__o21a_1 _28001_ (.A1(_11187_),
    .A2(_11202_),
    .B1(_11326_),
    .X(_11327_));
 sky130_fd_sc_hd__nand2_1 _28002_ (.A(_11144_),
    .B(_11128_),
    .Y(_11328_));
 sky130_fd_sc_hd__o21a_2 _28003_ (.A1(_11126_),
    .A2(_11145_),
    .B1(_11328_),
    .X(_11329_));
 sky130_fd_sc_hd__buf_2 _28004_ (.A(_11050_),
    .X(_11330_));
 sky130_fd_sc_hd__or2_1 _28005_ (.A(_11195_),
    .B(_11199_),
    .X(_11331_));
 sky130_fd_sc_hd__o21a_2 _28006_ (.A1(_11194_),
    .A2(_11200_),
    .B1(_11331_),
    .X(_11332_));
 sky130_vsdinv _28007_ (.A(_11057_),
    .Y(_11333_));
 sky130_fd_sc_hd__nor2_1 _28008_ (.A(_11196_),
    .B(_11197_),
    .Y(_11334_));
 sky130_fd_sc_hd__o21ba_4 _28009_ (.A1(_11333_),
    .A2(_11198_),
    .B1_N(_11334_),
    .X(_11335_));
 sky130_fd_sc_hd__o21a_2 _28010_ (.A1(_07820_),
    .A2(_08721_),
    .B1(_09283_),
    .X(_11336_));
 sky130_fd_sc_hd__nand3_4 _28011_ (.A(_09283_),
    .B(_07820_),
    .C(_05815_),
    .Y(_11337_));
 sky130_fd_sc_hd__nand2_2 _28012_ (.A(_11336_),
    .B(_11337_),
    .Y(_11338_));
 sky130_fd_sc_hd__xor2_4 _28013_ (.A(_11333_),
    .B(_11338_),
    .X(_11339_));
 sky130_fd_sc_hd__a21bo_2 _28014_ (.A1(_11141_),
    .A2(_11139_),
    .B1_N(_11140_),
    .X(_11340_));
 sky130_fd_sc_hd__xnor2_4 _28015_ (.A(_11339_),
    .B(_11340_),
    .Y(_11341_));
 sky130_fd_sc_hd__xnor2_4 _28016_ (.A(_11335_),
    .B(_11341_),
    .Y(_11342_));
 sky130_fd_sc_hd__xnor2_4 _28017_ (.A(_11332_),
    .B(_11342_),
    .Y(_11343_));
 sky130_fd_sc_hd__xor2_4 _28018_ (.A(net415),
    .B(_11343_),
    .X(_11344_));
 sky130_fd_sc_hd__xor2_4 _28019_ (.A(_11329_),
    .B(_11344_),
    .X(_11345_));
 sky130_fd_sc_hd__xnor2_2 _28020_ (.A(_11327_),
    .B(_11345_),
    .Y(_11346_));
 sky130_fd_sc_hd__a21o_1 _28021_ (.A1(_11324_),
    .A2(_11325_),
    .B1(_11346_),
    .X(_11347_));
 sky130_fd_sc_hd__nand3b_4 _28022_ (.A_N(_11323_),
    .B(_11346_),
    .C(_11325_),
    .Y(_11348_));
 sky130_vsdinv _28023_ (.A(_11205_),
    .Y(_11349_));
 sky130_fd_sc_hd__o21ai_2 _28024_ (.A1(_11349_),
    .A2(_11184_),
    .B1(_11186_),
    .Y(_11350_));
 sky130_fd_sc_hd__a21o_1 _28025_ (.A1(_11347_),
    .A2(_11348_),
    .B1(_11350_),
    .X(_11351_));
 sky130_fd_sc_hd__nand3_4 _28026_ (.A(_11347_),
    .B(_11350_),
    .C(_11348_),
    .Y(_11352_));
 sky130_fd_sc_hd__nor2_8 _28027_ (.A(_11079_),
    .B(_11215_),
    .Y(_11353_));
 sky130_fd_sc_hd__a21oi_4 _28028_ (.A1(_09978_),
    .A2(_11218_),
    .B1(_11353_),
    .Y(_11354_));
 sky130_fd_sc_hd__nor3b_2 _28029_ (.A(_10609_),
    .B(_10764_),
    .C_N(_11215_),
    .Y(_11355_));
 sky130_vsdinv _28030_ (.A(_11355_),
    .Y(_11356_));
 sky130_fd_sc_hd__o211a_1 _28031_ (.A1(_11079_),
    .A2(_11215_),
    .B1(_11356_),
    .C1(_09791_),
    .X(_11357_));
 sky130_vsdinv _28032_ (.A(_11353_),
    .Y(_11358_));
 sky130_fd_sc_hd__a21o_1 _28033_ (.A1(_11358_),
    .A2(_11356_),
    .B1(_09791_),
    .X(_11359_));
 sky130_fd_sc_hd__and2b_1 _28034_ (.A_N(_11357_),
    .B(_11359_),
    .X(_11360_));
 sky130_fd_sc_hd__buf_6 _28035_ (.A(_11360_),
    .X(_11361_));
 sky130_vsdinv _28036_ (.A(_11361_),
    .Y(_11362_));
 sky130_fd_sc_hd__buf_4 _28037_ (.A(_11362_),
    .X(_11363_));
 sky130_fd_sc_hd__nand2_1 _28038_ (.A(_11203_),
    .B(_11191_),
    .Y(_11364_));
 sky130_fd_sc_hd__o21ai_2 _28039_ (.A1(_11189_),
    .A2(_11204_),
    .B1(_11364_),
    .Y(_11365_));
 sky130_fd_sc_hd__xor2_2 _28040_ (.A(_11363_),
    .B(_11365_),
    .X(_11366_));
 sky130_fd_sc_hd__xnor2_1 _28041_ (.A(_11354_),
    .B(_11366_),
    .Y(_11367_));
 sky130_fd_sc_hd__a21bo_1 _28042_ (.A1(_11351_),
    .A2(_11352_),
    .B1_N(_11367_),
    .X(_11368_));
 sky130_fd_sc_hd__nand3b_4 _28043_ (.A_N(_11367_),
    .B(_11351_),
    .C(_11352_),
    .Y(_11369_));
 sky130_fd_sc_hd__a21oi_1 _28044_ (.A1(_11211_),
    .A2(_11207_),
    .B1(_11209_),
    .Y(_11370_));
 sky130_fd_sc_hd__o21ai_2 _28045_ (.A1(_11223_),
    .A2(_11370_),
    .B1(_11212_),
    .Y(_11371_));
 sky130_fd_sc_hd__a21o_2 _28046_ (.A1(_11368_),
    .A2(_11369_),
    .B1(_11371_),
    .X(_11372_));
 sky130_fd_sc_hd__nand3_4 _28047_ (.A(_11371_),
    .B(_11368_),
    .C(_11369_),
    .Y(_11373_));
 sky130_fd_sc_hd__and2_1 _28048_ (.A(_11221_),
    .B(_11219_),
    .X(_11374_));
 sky130_fd_sc_hd__o21bai_4 _28049_ (.A1(_11214_),
    .A2(_11222_),
    .B1_N(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__xor2_4 _28050_ (.A(_10178_),
    .B(_11375_),
    .X(_11376_));
 sky130_fd_sc_hd__a21oi_2 _28051_ (.A1(_11372_),
    .A2(_11373_),
    .B1(_11376_),
    .Y(_11377_));
 sky130_fd_sc_hd__nand3_4 _28052_ (.A(_11372_),
    .B(_11376_),
    .C(_11373_),
    .Y(_11378_));
 sky130_vsdinv _28053_ (.A(_11231_),
    .Y(_11379_));
 sky130_fd_sc_hd__o21ai_2 _28054_ (.A1(_11379_),
    .A2(_11227_),
    .B1(_11228_),
    .Y(_11380_));
 sky130_fd_sc_hd__nand3b_4 _28055_ (.A_N(_11377_),
    .B(_11378_),
    .C(_11380_),
    .Y(_11381_));
 sky130_vsdinv _28056_ (.A(_11378_),
    .Y(_11382_));
 sky130_fd_sc_hd__o21bai_2 _28057_ (.A1(_11377_),
    .A2(_11382_),
    .B1_N(_11380_),
    .Y(_11383_));
 sky130_fd_sc_hd__o2bb2ai_2 _28058_ (.A1_N(_11381_),
    .A2_N(_11383_),
    .B1(_11243_),
    .B2(_11230_),
    .Y(_11384_));
 sky130_fd_sc_hd__a21oi_4 _28059_ (.A1(_11091_),
    .A2(_11086_),
    .B1(_10812_),
    .Y(_11385_));
 sky130_fd_sc_hd__nand3_4 _28060_ (.A(_11383_),
    .B(_11381_),
    .C(_11385_),
    .Y(_11386_));
 sky130_vsdinv _28061_ (.A(_11245_),
    .Y(_11387_));
 sky130_fd_sc_hd__a21oi_2 _28062_ (.A1(_11232_),
    .A2(_11236_),
    .B1(_11237_),
    .Y(_11388_));
 sky130_fd_sc_hd__o21ai_4 _28063_ (.A1(_11387_),
    .A2(_11388_),
    .B1(_11238_),
    .Y(_11389_));
 sky130_fd_sc_hd__a21o_1 _28064_ (.A1(_11384_),
    .A2(_11386_),
    .B1(_11389_),
    .X(_11390_));
 sky130_fd_sc_hd__nand3_4 _28065_ (.A(_11384_),
    .B(_11389_),
    .C(_11386_),
    .Y(_11391_));
 sky130_fd_sc_hd__nand2_2 _28066_ (.A(_11390_),
    .B(_11391_),
    .Y(_11392_));
 sky130_fd_sc_hd__a21boi_1 _28067_ (.A1(_11269_),
    .A2(_11249_),
    .B1_N(_11250_),
    .Y(_11393_));
 sky130_fd_sc_hd__xor2_1 _28068_ (.A(_11392_),
    .B(_11393_),
    .X(_02668_));
 sky130_fd_sc_hd__or2_1 _28069_ (.A(_11332_),
    .B(_11342_),
    .X(_11394_));
 sky130_fd_sc_hd__o21a_1 _28070_ (.A1(_11187_),
    .A2(_11343_),
    .B1(_11394_),
    .X(_11395_));
 sky130_vsdinv _28071_ (.A(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__nand2_1 _28072_ (.A(_11288_),
    .B(_11275_),
    .Y(_11397_));
 sky130_fd_sc_hd__o21a_1 _28073_ (.A1(_11273_),
    .A2(_11289_),
    .B1(_11397_),
    .X(_11398_));
 sky130_fd_sc_hd__and2_1 _28074_ (.A(_11340_),
    .B(_11339_),
    .X(_11399_));
 sky130_fd_sc_hd__o21bai_4 _28075_ (.A1(_11335_),
    .A2(_11341_),
    .B1_N(_11399_),
    .Y(_11400_));
 sky130_fd_sc_hd__a21boi_4 _28076_ (.A1(_11336_),
    .A2(_11057_),
    .B1_N(_11337_),
    .Y(_11401_));
 sky130_fd_sc_hd__a21bo_2 _28077_ (.A1(_11285_),
    .A2(_11283_),
    .B1_N(_11284_),
    .X(_11402_));
 sky130_fd_sc_hd__xnor2_4 _28078_ (.A(_11339_),
    .B(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__xor2_4 _28079_ (.A(_11401_),
    .B(_11403_),
    .X(_11404_));
 sky130_fd_sc_hd__xnor2_4 _28080_ (.A(_11400_),
    .B(_11404_),
    .Y(_11405_));
 sky130_fd_sc_hd__xor2_4 _28081_ (.A(net415),
    .B(_11405_),
    .X(_11406_));
 sky130_fd_sc_hd__xor2_2 _28082_ (.A(_11398_),
    .B(_11406_),
    .X(_11407_));
 sky130_fd_sc_hd__xor2_1 _28083_ (.A(_11396_),
    .B(_11407_),
    .X(_11408_));
 sky130_vsdinv _28084_ (.A(_11408_),
    .Y(_11409_));
 sky130_fd_sc_hd__nand2_1 _28085_ (.A(_11320_),
    .B(_11293_),
    .Y(_11410_));
 sky130_fd_sc_hd__o21a_1 _28086_ (.A1(_11291_),
    .A2(_11321_),
    .B1(_11410_),
    .X(_11411_));
 sky130_fd_sc_hd__nor2_1 _28087_ (.A(_11276_),
    .B(_11281_),
    .Y(_11412_));
 sky130_fd_sc_hd__o21ba_1 _28088_ (.A1(_11282_),
    .A2(_11287_),
    .B1_N(_11412_),
    .X(_11413_));
 sky130_fd_sc_hd__nor2_1 _28089_ (.A(_11295_),
    .B(_11300_),
    .Y(_11414_));
 sky130_fd_sc_hd__o21bai_2 _28090_ (.A1(_11294_),
    .A2(_11301_),
    .B1_N(_11414_),
    .Y(_11415_));
 sky130_fd_sc_hd__a2bb2oi_4 _28091_ (.A1_N(_14299_),
    .A2_N(_11278_),
    .B1(_11277_),
    .B2(_11279_),
    .Y(_11416_));
 sky130_fd_sc_hd__and2_2 _28092_ (.A(_09388_),
    .B(_08157_),
    .X(_11417_));
 sky130_fd_sc_hd__nand3_4 _28093_ (.A(_11132_),
    .B(_11133_),
    .C(_07769_),
    .Y(_11418_));
 sky130_fd_sc_hd__a22o_2 _28094_ (.A1(_10515_),
    .A2(_08070_),
    .B1(_10516_),
    .B2(_07778_),
    .X(_11419_));
 sky130_fd_sc_hd__o21ai_4 _28095_ (.A1(_14292_),
    .A2(_11418_),
    .B1(_11419_),
    .Y(_11420_));
 sky130_fd_sc_hd__xor2_4 _28096_ (.A(_11417_),
    .B(_11420_),
    .X(_11421_));
 sky130_fd_sc_hd__xnor2_2 _28097_ (.A(_11416_),
    .B(_11421_),
    .Y(_11422_));
 sky130_fd_sc_hd__and2_1 _28098_ (.A(_12778_),
    .B(_06059_),
    .X(_11423_));
 sky130_fd_sc_hd__buf_4 _28099_ (.A(_11423_),
    .X(_11424_));
 sky130_fd_sc_hd__or4_4 _28100_ (.A(_14011_),
    .B(_14016_),
    .C(_14275_),
    .D(_14279_),
    .X(_11425_));
 sky130_fd_sc_hd__a22o_1 _28101_ (.A1(_08857_),
    .A2(_08480_),
    .B1(_08423_),
    .B2(_08492_),
    .X(_11426_));
 sky130_fd_sc_hd__nand2_4 _28102_ (.A(_11425_),
    .B(_11426_),
    .Y(_11427_));
 sky130_fd_sc_hd__xor2_4 _28103_ (.A(_11424_),
    .B(_11427_),
    .X(_11428_));
 sky130_fd_sc_hd__xor2_2 _28104_ (.A(_11422_),
    .B(_11428_),
    .X(_11429_));
 sky130_fd_sc_hd__xnor2_1 _28105_ (.A(_11415_),
    .B(_11429_),
    .Y(_11430_));
 sky130_fd_sc_hd__xor2_1 _28106_ (.A(_11413_),
    .B(_11430_),
    .X(_11431_));
 sky130_vsdinv _28107_ (.A(_11431_),
    .Y(_11432_));
 sky130_fd_sc_hd__and2_1 _28108_ (.A(_11318_),
    .B(_11304_),
    .X(_11433_));
 sky130_fd_sc_hd__o21bai_4 _28109_ (.A1(_11302_),
    .A2(_11319_),
    .B1_N(_11433_),
    .Y(_11434_));
 sky130_fd_sc_hd__a2bb2oi_4 _28110_ (.A1_N(_14316_),
    .A2_N(_11297_),
    .B1(_11296_),
    .B2(_11298_),
    .Y(_11435_));
 sky130_fd_sc_hd__a2bb2oi_4 _28111_ (.A1_N(_14335_),
    .A2_N(_11306_),
    .B1(_11305_),
    .B2(_11307_),
    .Y(_11436_));
 sky130_fd_sc_hd__nand2_2 _28112_ (.A(net437),
    .B(_07570_),
    .Y(_11437_));
 sky130_fd_sc_hd__or4_4 _28113_ (.A(_13986_),
    .B(_13991_),
    .C(_14309_),
    .D(_14314_),
    .X(_11438_));
 sky130_fd_sc_hd__a22o_1 _28114_ (.A1(_10672_),
    .A2(_07473_),
    .B1(_11009_),
    .B2(_08885_),
    .X(_11439_));
 sky130_fd_sc_hd__nand2_2 _28115_ (.A(_11438_),
    .B(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__xnor2_4 _28116_ (.A(_11437_),
    .B(_11440_),
    .Y(_11441_));
 sky130_fd_sc_hd__xnor2_4 _28117_ (.A(_11436_),
    .B(_11441_),
    .Y(_11442_));
 sky130_fd_sc_hd__xnor2_4 _28118_ (.A(_11435_),
    .B(_11442_),
    .Y(_11443_));
 sky130_fd_sc_hd__or2b_2 _28119_ (.A(_11316_),
    .B_N(_11311_),
    .X(_11444_));
 sky130_fd_sc_hd__o21ai_4 _28120_ (.A1(_11309_),
    .A2(_11317_),
    .B1(_11444_),
    .Y(_11445_));
 sky130_fd_sc_hd__and2_2 _28121_ (.A(_11162_),
    .B(_07028_),
    .X(_11446_));
 sky130_fd_sc_hd__nand3_4 _28122_ (.A(_13973_),
    .B(_11166_),
    .C(_06762_),
    .Y(_11447_));
 sky130_fd_sc_hd__a22o_2 _28123_ (.A1(_11018_),
    .A2(_06762_),
    .B1(_13979_),
    .B2(_06941_),
    .X(_11448_));
 sky130_fd_sc_hd__o21ai_4 _28124_ (.A1(_08332_),
    .A2(_11447_),
    .B1(_11448_),
    .Y(_11449_));
 sky130_fd_sc_hd__xor2_4 _28125_ (.A(_11446_),
    .B(_11449_),
    .X(_11450_));
 sky130_fd_sc_hd__nand3b_2 _28126_ (.A_N(_11313_),
    .B(_11025_),
    .C(_14360_),
    .Y(_11451_));
 sky130_fd_sc_hd__o31ai_4 _28127_ (.A1(_13968_),
    .A2(_14348_),
    .A3(_11315_),
    .B1(_11451_),
    .Y(_11452_));
 sky130_fd_sc_hd__and2_2 _28128_ (.A(_11028_),
    .B(_07747_),
    .X(_11453_));
 sky130_fd_sc_hd__nand2_2 _28129_ (.A(_13962_),
    .B(_06431_),
    .Y(_11454_));
 sky130_fd_sc_hd__and2b_1 _28130_ (.A_N(_06288_),
    .B(_09025_),
    .X(_11455_));
 sky130_fd_sc_hd__xor2_4 _28131_ (.A(_11454_),
    .B(_11455_),
    .X(_11456_));
 sky130_fd_sc_hd__xor2_4 _28132_ (.A(_11453_),
    .B(_11456_),
    .X(_11457_));
 sky130_fd_sc_hd__xor2_4 _28133_ (.A(_11452_),
    .B(_11457_),
    .X(_11458_));
 sky130_fd_sc_hd__xor2_4 _28134_ (.A(_11450_),
    .B(_11458_),
    .X(_11459_));
 sky130_fd_sc_hd__xnor2_4 _28135_ (.A(_11445_),
    .B(_11459_),
    .Y(_11460_));
 sky130_fd_sc_hd__xor2_4 _28136_ (.A(_11443_),
    .B(_11460_),
    .X(_11461_));
 sky130_fd_sc_hd__xnor2_4 _28137_ (.A(_11434_),
    .B(_11461_),
    .Y(_11462_));
 sky130_fd_sc_hd__xor2_4 _28138_ (.A(_11432_),
    .B(_11462_),
    .X(_11463_));
 sky130_fd_sc_hd__xor2_2 _28139_ (.A(_11411_),
    .B(_11463_),
    .X(_11464_));
 sky130_fd_sc_hd__nor2_1 _28140_ (.A(_11409_),
    .B(_11464_),
    .Y(_11465_));
 sky130_vsdinv _28141_ (.A(_11465_),
    .Y(_11466_));
 sky130_fd_sc_hd__nand2_2 _28142_ (.A(_11464_),
    .B(_11409_),
    .Y(_11467_));
 sky130_fd_sc_hd__a21o_1 _28143_ (.A1(_11325_),
    .A2(_11346_),
    .B1(_11323_),
    .X(_11468_));
 sky130_fd_sc_hd__a21oi_1 _28144_ (.A1(_11466_),
    .A2(_11467_),
    .B1(_11468_),
    .Y(_11469_));
 sky130_vsdinv _28145_ (.A(_11469_),
    .Y(_11470_));
 sky130_fd_sc_hd__nand3b_4 _28146_ (.A_N(_11465_),
    .B(_11467_),
    .C(_11468_),
    .Y(_11471_));
 sky130_fd_sc_hd__a21oi_4 _28147_ (.A1(_09978_),
    .A2(_11356_),
    .B1(_11353_),
    .Y(_11472_));
 sky130_fd_sc_hd__clkbuf_8 _28148_ (.A(_11472_),
    .X(_11473_));
 sky130_fd_sc_hd__or2b_2 _28149_ (.A(_11327_),
    .B_N(_11345_),
    .X(_11474_));
 sky130_fd_sc_hd__or2_2 _28150_ (.A(_11329_),
    .B(_11344_),
    .X(_11475_));
 sky130_fd_sc_hd__clkbuf_4 _28151_ (.A(_11362_),
    .X(_11476_));
 sky130_fd_sc_hd__a21o_1 _28152_ (.A1(_11474_),
    .A2(_11475_),
    .B1(_11476_),
    .X(_11477_));
 sky130_fd_sc_hd__nand3_4 _28153_ (.A(_11474_),
    .B(_11476_),
    .C(_11475_),
    .Y(_11478_));
 sky130_fd_sc_hd__nand2_2 _28154_ (.A(_11477_),
    .B(_11478_),
    .Y(_11479_));
 sky130_fd_sc_hd__xor2_4 _28155_ (.A(_11473_),
    .B(_11479_),
    .X(_11480_));
 sky130_fd_sc_hd__a21oi_2 _28156_ (.A1(_11470_),
    .A2(_11471_),
    .B1(_11480_),
    .Y(_11481_));
 sky130_fd_sc_hd__nand3b_4 _28157_ (.A_N(_11469_),
    .B(_11480_),
    .C(_11471_),
    .Y(_11482_));
 sky130_vsdinv _28158_ (.A(_11482_),
    .Y(_11483_));
 sky130_fd_sc_hd__nand2_2 _28159_ (.A(_11369_),
    .B(_11352_),
    .Y(_11484_));
 sky130_fd_sc_hd__o21bai_4 _28160_ (.A1(_11481_),
    .A2(_11483_),
    .B1_N(_11484_),
    .Y(_11485_));
 sky130_fd_sc_hd__a21o_1 _28161_ (.A1(_11470_),
    .A2(_11471_),
    .B1(_11480_),
    .X(_11486_));
 sky130_fd_sc_hd__nand3_4 _28162_ (.A(_11486_),
    .B(_11482_),
    .C(_11484_),
    .Y(_11487_));
 sky130_fd_sc_hd__or2_1 _28163_ (.A(_11189_),
    .B(_11204_),
    .X(_11488_));
 sky130_fd_sc_hd__buf_4 _28164_ (.A(_11476_),
    .X(_11489_));
 sky130_fd_sc_hd__a21o_1 _28165_ (.A1(_11488_),
    .A2(_11364_),
    .B1(_11489_),
    .X(_11490_));
 sky130_fd_sc_hd__o21a_4 _28166_ (.A1(_11354_),
    .A2(_11366_),
    .B1(_11490_),
    .X(_11491_));
 sky130_fd_sc_hd__xor2_4 _28167_ (.A(net413),
    .B(_11491_),
    .X(_11492_));
 sky130_fd_sc_hd__a21oi_4 _28168_ (.A1(_11485_),
    .A2(_11487_),
    .B1(_11492_),
    .Y(_11493_));
 sky130_fd_sc_hd__nand3_4 _28169_ (.A(_11485_),
    .B(_11492_),
    .C(_11487_),
    .Y(_11494_));
 sky130_vsdinv _28170_ (.A(_11494_),
    .Y(_11495_));
 sky130_fd_sc_hd__a21boi_4 _28171_ (.A1(_11372_),
    .A2(_11376_),
    .B1_N(_11373_),
    .Y(_11496_));
 sky130_fd_sc_hd__o21ai_4 _28172_ (.A1(_11493_),
    .A2(_11495_),
    .B1(_11496_),
    .Y(_11497_));
 sky130_fd_sc_hd__nand2_1 _28173_ (.A(_11378_),
    .B(_11373_),
    .Y(_11498_));
 sky130_fd_sc_hd__nand3b_4 _28174_ (.A_N(_11493_),
    .B(_11494_),
    .C(_11498_),
    .Y(_11499_));
 sky130_fd_sc_hd__and2_2 _28175_ (.A(_11375_),
    .B(_10178_),
    .X(_11500_));
 sky130_fd_sc_hd__a21o_1 _28176_ (.A1(_11497_),
    .A2(_11499_),
    .B1(_11500_),
    .X(_11501_));
 sky130_fd_sc_hd__nand3_4 _28177_ (.A(_11497_),
    .B(_11499_),
    .C(_11500_),
    .Y(_11502_));
 sky130_fd_sc_hd__nand2_2 _28178_ (.A(_11386_),
    .B(_11381_),
    .Y(_11503_));
 sky130_fd_sc_hd__a21oi_4 _28179_ (.A1(_11501_),
    .A2(_11502_),
    .B1(_11503_),
    .Y(_11504_));
 sky130_fd_sc_hd__nand3_2 _28180_ (.A(_11501_),
    .B(_11503_),
    .C(_11502_),
    .Y(_11505_));
 sky130_vsdinv _28181_ (.A(_11505_),
    .Y(_11506_));
 sky130_fd_sc_hd__nor2_8 _28182_ (.A(_11504_),
    .B(_11506_),
    .Y(_11507_));
 sky130_fd_sc_hd__nor2_4 _28183_ (.A(_11392_),
    .B(_11251_),
    .Y(_11508_));
 sky130_fd_sc_hd__a21oi_2 _28184_ (.A1(_11384_),
    .A2(_11386_),
    .B1(_11389_),
    .Y(_11509_));
 sky130_fd_sc_hd__a21oi_4 _28185_ (.A1(_11250_),
    .A2(_11391_),
    .B1(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__a21oi_2 _28186_ (.A1(_11269_),
    .A2(_11508_),
    .B1(_11510_),
    .Y(_11511_));
 sky130_fd_sc_hd__xnor2_1 _28187_ (.A(_11507_),
    .B(_11511_),
    .Y(_02669_));
 sky130_fd_sc_hd__nand2_2 _28188_ (.A(_11407_),
    .B(_11396_),
    .Y(_11512_));
 sky130_fd_sc_hd__or2_2 _28189_ (.A(_11398_),
    .B(_11406_),
    .X(_11513_));
 sky130_fd_sc_hd__a21o_1 _28190_ (.A1(_11512_),
    .A2(_11513_),
    .B1(_11362_),
    .X(_11514_));
 sky130_fd_sc_hd__nand3_4 _28191_ (.A(_11512_),
    .B(_11363_),
    .C(_11513_),
    .Y(_11515_));
 sky130_fd_sc_hd__nand2_1 _28192_ (.A(_11514_),
    .B(_11515_),
    .Y(_11516_));
 sky130_fd_sc_hd__xor2_1 _28193_ (.A(_11472_),
    .B(_11516_),
    .X(_11517_));
 sky130_vsdinv _28194_ (.A(_11517_),
    .Y(_11518_));
 sky130_fd_sc_hd__and2b_1 _28195_ (.A_N(_11463_),
    .B(_11411_),
    .X(_11519_));
 sky130_fd_sc_hd__or2b_1 _28196_ (.A(_11411_),
    .B_N(_11463_),
    .X(_11520_));
 sky130_fd_sc_hd__o21a_1 _28197_ (.A1(_11409_),
    .A2(_11519_),
    .B1(_11520_),
    .X(_11521_));
 sky130_fd_sc_hd__nand2_1 _28198_ (.A(_11404_),
    .B(_11400_),
    .Y(_11522_));
 sky130_fd_sc_hd__o21a_1 _28199_ (.A1(_11051_),
    .A2(_11405_),
    .B1(_11522_),
    .X(_11523_));
 sky130_vsdinv _28200_ (.A(_11523_),
    .Y(_11524_));
 sky130_fd_sc_hd__nand2_1 _28201_ (.A(_11429_),
    .B(_11415_),
    .Y(_11525_));
 sky130_fd_sc_hd__o21a_1 _28202_ (.A1(_11413_),
    .A2(_11430_),
    .B1(_11525_),
    .X(_11526_));
 sky130_fd_sc_hd__and2_1 _28203_ (.A(_11402_),
    .B(_11339_),
    .X(_11527_));
 sky130_fd_sc_hd__o21bai_4 _28204_ (.A1(_11401_),
    .A2(_11403_),
    .B1_N(_11527_),
    .Y(_11528_));
 sky130_fd_sc_hd__clkinv_4 _28205_ (.A(_11424_),
    .Y(_11529_));
 sky130_fd_sc_hd__o21ai_4 _28206_ (.A1(_11529_),
    .A2(_11427_),
    .B1(_11425_),
    .Y(_11530_));
 sky130_fd_sc_hd__xnor2_4 _28207_ (.A(_11339_),
    .B(_11530_),
    .Y(_11531_));
 sky130_fd_sc_hd__xor2_4 _28208_ (.A(_11401_),
    .B(_11531_),
    .X(_11532_));
 sky130_fd_sc_hd__xnor2_4 _28209_ (.A(_11528_),
    .B(_11532_),
    .Y(_11533_));
 sky130_fd_sc_hd__xor2_4 _28210_ (.A(net415),
    .B(_11533_),
    .X(_11534_));
 sky130_fd_sc_hd__xor2_2 _28211_ (.A(_11526_),
    .B(_11534_),
    .X(_11535_));
 sky130_fd_sc_hd__xor2_1 _28212_ (.A(_11524_),
    .B(_11535_),
    .X(_11536_));
 sky130_vsdinv _28213_ (.A(_11536_),
    .Y(_11537_));
 sky130_fd_sc_hd__and2_1 _28214_ (.A(_11461_),
    .B(_11434_),
    .X(_11538_));
 sky130_fd_sc_hd__o21ba_2 _28215_ (.A1(_11432_),
    .A2(_11462_),
    .B1_N(_11538_),
    .X(_11539_));
 sky130_fd_sc_hd__nor2_1 _28216_ (.A(_11416_),
    .B(_11421_),
    .Y(_11540_));
 sky130_fd_sc_hd__o21ba_1 _28217_ (.A1(_11422_),
    .A2(_11428_),
    .B1_N(_11540_),
    .X(_11541_));
 sky130_fd_sc_hd__nand2_2 _28218_ (.A(_10984_),
    .B(_08596_),
    .Y(_11542_));
 sky130_fd_sc_hd__nand2_8 _28219_ (.A(_12778_),
    .B(_09379_),
    .Y(_11543_));
 sky130_fd_sc_hd__xnor2_4 _28220_ (.A(_11542_),
    .B(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__xor2_4 _28221_ (.A(_11424_),
    .B(_11544_),
    .X(_11545_));
 sky130_fd_sc_hd__a2bb2oi_4 _28222_ (.A1_N(_14293_),
    .A2_N(_11418_),
    .B1(_11417_),
    .B2(_11419_),
    .Y(_11546_));
 sky130_fd_sc_hd__and2_2 _28223_ (.A(_06472_),
    .B(_08480_),
    .X(_11547_));
 sky130_fd_sc_hd__nand3_4 _28224_ (.A(_10991_),
    .B(_11133_),
    .C(_08064_),
    .Y(_11548_));
 sky130_fd_sc_hd__a22o_2 _28225_ (.A1(_10515_),
    .A2(_07778_),
    .B1(_11133_),
    .B2(_08488_),
    .X(_11549_));
 sky130_fd_sc_hd__o21ai_4 _28226_ (.A1(_14286_),
    .A2(_11548_),
    .B1(_11549_),
    .Y(_11550_));
 sky130_fd_sc_hd__xor2_4 _28227_ (.A(_11547_),
    .B(_11550_),
    .X(_11551_));
 sky130_fd_sc_hd__xnor2_2 _28228_ (.A(_11546_),
    .B(_11551_),
    .Y(_11552_));
 sky130_fd_sc_hd__xor2_2 _28229_ (.A(_11545_),
    .B(_11552_),
    .X(_11553_));
 sky130_fd_sc_hd__nor2_1 _28230_ (.A(_11436_),
    .B(_11441_),
    .Y(_11554_));
 sky130_fd_sc_hd__o21bai_2 _28231_ (.A1(_11435_),
    .A2(_11442_),
    .B1_N(_11554_),
    .Y(_11555_));
 sky130_fd_sc_hd__xnor2_1 _28232_ (.A(_11553_),
    .B(_11555_),
    .Y(_11556_));
 sky130_fd_sc_hd__xor2_1 _28233_ (.A(_11541_),
    .B(_11556_),
    .X(_11557_));
 sky130_vsdinv _28234_ (.A(_11557_),
    .Y(_11558_));
 sky130_fd_sc_hd__and2_1 _28235_ (.A(_11459_),
    .B(_11445_),
    .X(_11559_));
 sky130_fd_sc_hd__o21bai_4 _28236_ (.A1(_11443_),
    .A2(_11460_),
    .B1_N(_11559_),
    .Y(_11560_));
 sky130_fd_sc_hd__o21a_2 _28237_ (.A1(_11437_),
    .A2(_11440_),
    .B1(_11438_),
    .X(_11561_));
 sky130_fd_sc_hd__a2bb2oi_4 _28238_ (.A1_N(_14329_),
    .A2_N(_11447_),
    .B1(_11446_),
    .B2(_11448_),
    .Y(_11562_));
 sky130_fd_sc_hd__nand2_2 _28239_ (.A(net437),
    .B(_10829_),
    .Y(_11563_));
 sky130_fd_sc_hd__or4_4 _28240_ (.A(_13985_),
    .B(_13991_),
    .C(_14304_),
    .D(_14308_),
    .X(_11564_));
 sky130_fd_sc_hd__a22o_1 _28241_ (.A1(_10672_),
    .A2(_07467_),
    .B1(_07103_),
    .B2(_07569_),
    .X(_11565_));
 sky130_fd_sc_hd__nand2_2 _28242_ (.A(_11564_),
    .B(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__xnor2_4 _28243_ (.A(_11563_),
    .B(_11566_),
    .Y(_11567_));
 sky130_fd_sc_hd__xnor2_4 _28244_ (.A(_11562_),
    .B(_11567_),
    .Y(_11568_));
 sky130_fd_sc_hd__xnor2_4 _28245_ (.A(_11561_),
    .B(_11568_),
    .Y(_11569_));
 sky130_fd_sc_hd__or2b_2 _28246_ (.A(_11457_),
    .B_N(_11452_),
    .X(_11570_));
 sky130_fd_sc_hd__o21ai_4 _28247_ (.A1(_11450_),
    .A2(_11458_),
    .B1(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__and2_2 _28248_ (.A(_11162_),
    .B(_07199_),
    .X(_11572_));
 sky130_fd_sc_hd__nand3_4 _28249_ (.A(_13973_),
    .B(_11166_),
    .C(_06941_),
    .Y(_11573_));
 sky130_fd_sc_hd__a22o_2 _28250_ (.A1(_08397_),
    .A2(_06941_),
    .B1(_13979_),
    .B2(_07028_),
    .X(_11574_));
 sky130_fd_sc_hd__o21ai_4 _28251_ (.A1(_14321_),
    .A2(_11573_),
    .B1(_11574_),
    .Y(_11575_));
 sky130_fd_sc_hd__xor2_4 _28252_ (.A(_11572_),
    .B(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__nand3b_4 _28253_ (.A_N(_11454_),
    .B(_11025_),
    .C(_08338_),
    .Y(_11577_));
 sky130_fd_sc_hd__o31ai_4 _28254_ (.A1(_11024_),
    .A2(_14341_),
    .A3(_11456_),
    .B1(_11577_),
    .Y(_11578_));
 sky130_fd_sc_hd__and2_2 _28255_ (.A(_11028_),
    .B(_06761_),
    .X(_11579_));
 sky130_fd_sc_hd__nand2_2 _28256_ (.A(_11030_),
    .B(_07746_),
    .Y(_11580_));
 sky130_fd_sc_hd__and2b_2 _28257_ (.A_N(_06165_),
    .B(_12805_),
    .X(_11581_));
 sky130_fd_sc_hd__xor2_4 _28258_ (.A(_11580_),
    .B(_11581_),
    .X(_11582_));
 sky130_fd_sc_hd__xor2_4 _28259_ (.A(_11579_),
    .B(_11582_),
    .X(_11583_));
 sky130_fd_sc_hd__xor2_4 _28260_ (.A(_11578_),
    .B(_11583_),
    .X(_11584_));
 sky130_fd_sc_hd__xor2_4 _28261_ (.A(_11576_),
    .B(_11584_),
    .X(_11585_));
 sky130_fd_sc_hd__xnor2_4 _28262_ (.A(_11571_),
    .B(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__xor2_4 _28263_ (.A(_11569_),
    .B(_11586_),
    .X(_11587_));
 sky130_fd_sc_hd__xnor2_4 _28264_ (.A(_11560_),
    .B(_11587_),
    .Y(_11588_));
 sky130_fd_sc_hd__xor2_4 _28265_ (.A(_11558_),
    .B(_11588_),
    .X(_11589_));
 sky130_fd_sc_hd__xor2_4 _28266_ (.A(_11539_),
    .B(_11589_),
    .X(_11590_));
 sky130_fd_sc_hd__nor2_4 _28267_ (.A(_11537_),
    .B(_11590_),
    .Y(_11591_));
 sky130_fd_sc_hd__and2_1 _28268_ (.A(_11590_),
    .B(_11537_),
    .X(_11592_));
 sky130_fd_sc_hd__nor3_4 _28269_ (.A(_11521_),
    .B(_11591_),
    .C(_11592_),
    .Y(_11593_));
 sky130_fd_sc_hd__o21a_1 _28270_ (.A1(_11591_),
    .A2(_11592_),
    .B1(_11521_),
    .X(_11594_));
 sky130_fd_sc_hd__nor3_1 _28271_ (.A(_11518_),
    .B(_11593_),
    .C(_11594_),
    .Y(_11595_));
 sky130_vsdinv _28272_ (.A(_11595_),
    .Y(_11596_));
 sky130_fd_sc_hd__o21bai_2 _28273_ (.A1(_11593_),
    .A2(_11594_),
    .B1_N(_11517_),
    .Y(_11597_));
 sky130_fd_sc_hd__nand2_2 _28274_ (.A(_11482_),
    .B(_11471_),
    .Y(_11598_));
 sky130_fd_sc_hd__a21o_1 _28275_ (.A1(_11596_),
    .A2(_11597_),
    .B1(_11598_),
    .X(_11599_));
 sky130_fd_sc_hd__nand3_4 _28276_ (.A(_11598_),
    .B(_11596_),
    .C(_11597_),
    .Y(_11600_));
 sky130_vsdinv _28277_ (.A(_11472_),
    .Y(_11601_));
 sky130_fd_sc_hd__buf_6 _28278_ (.A(_11601_),
    .X(_11602_));
 sky130_fd_sc_hd__clkbuf_2 _28279_ (.A(_11602_),
    .X(_11603_));
 sky130_fd_sc_hd__a21boi_4 _28280_ (.A1(_11603_),
    .A2(_11478_),
    .B1_N(_11477_),
    .Y(_11604_));
 sky130_fd_sc_hd__xor2_4 _28281_ (.A(net413),
    .B(_11604_),
    .X(_11605_));
 sky130_fd_sc_hd__a21o_1 _28282_ (.A1(_11599_),
    .A2(_11600_),
    .B1(_11605_),
    .X(_11606_));
 sky130_vsdinv _28283_ (.A(_11492_),
    .Y(_11607_));
 sky130_fd_sc_hd__a21oi_1 _28284_ (.A1(_11486_),
    .A2(_11482_),
    .B1(_11484_),
    .Y(_11608_));
 sky130_fd_sc_hd__o21ai_2 _28285_ (.A1(_11607_),
    .A2(_11608_),
    .B1(_11487_),
    .Y(_11609_));
 sky130_fd_sc_hd__nand3_4 _28286_ (.A(_11599_),
    .B(_11605_),
    .C(_11600_),
    .Y(_11610_));
 sky130_fd_sc_hd__nand3_4 _28287_ (.A(_11606_),
    .B(_11609_),
    .C(_11610_),
    .Y(_11611_));
 sky130_fd_sc_hd__a21oi_2 _28288_ (.A1(_11599_),
    .A2(_11600_),
    .B1(_11605_),
    .Y(_11612_));
 sky130_vsdinv _28289_ (.A(_11610_),
    .Y(_11613_));
 sky130_fd_sc_hd__o21bai_4 _28290_ (.A1(_11612_),
    .A2(_11613_),
    .B1_N(_11609_),
    .Y(_11614_));
 sky130_fd_sc_hd__buf_4 _28291_ (.A(_11242_),
    .X(_11615_));
 sky130_fd_sc_hd__o2bb2ai_2 _28292_ (.A1_N(_11611_),
    .A2_N(_11614_),
    .B1(_11615_),
    .B2(_11491_),
    .Y(_11616_));
 sky130_fd_sc_hd__nor2_4 _28293_ (.A(_10813_),
    .B(_11491_),
    .Y(_11617_));
 sky130_fd_sc_hd__nand3_4 _28294_ (.A(_11614_),
    .B(_11617_),
    .C(_11611_),
    .Y(_11618_));
 sky130_fd_sc_hd__nor3_4 _28295_ (.A(_11496_),
    .B(_11493_),
    .C(_11495_),
    .Y(_11619_));
 sky130_fd_sc_hd__a21o_1 _28296_ (.A1(_11497_),
    .A2(_11500_),
    .B1(_11619_),
    .X(_11620_));
 sky130_fd_sc_hd__a21oi_4 _28297_ (.A1(_11616_),
    .A2(_11618_),
    .B1(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__a21oi_2 _28298_ (.A1(_11497_),
    .A2(_11500_),
    .B1(_11619_),
    .Y(_11622_));
 sky130_fd_sc_hd__a21oi_4 _28299_ (.A1(_11614_),
    .A2(_11611_),
    .B1(_11617_),
    .Y(_11623_));
 sky130_vsdinv _28300_ (.A(_11618_),
    .Y(_11624_));
 sky130_fd_sc_hd__nor3_4 _28301_ (.A(_11622_),
    .B(_11623_),
    .C(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__nor2_8 _28302_ (.A(_11621_),
    .B(_11625_),
    .Y(_11626_));
 sky130_fd_sc_hd__o21bai_1 _28303_ (.A1(_11504_),
    .A2(_11511_),
    .B1_N(_11506_),
    .Y(_11627_));
 sky130_fd_sc_hd__xor2_1 _28304_ (.A(_11626_),
    .B(_11627_),
    .X(_02670_));
 sky130_fd_sc_hd__or2_1 _28305_ (.A(_11546_),
    .B(_11551_),
    .X(_11628_));
 sky130_fd_sc_hd__o21a_2 _28306_ (.A1(_11545_),
    .A2(_11552_),
    .B1(_11628_),
    .X(_11629_));
 sky130_fd_sc_hd__nand2_2 _28307_ (.A(_09283_),
    .B(_08660_),
    .Y(_11630_));
 sky130_fd_sc_hd__xnor2_4 _28308_ (.A(_11543_),
    .B(_11630_),
    .Y(_11631_));
 sky130_fd_sc_hd__xor2_4 _28309_ (.A(_11529_),
    .B(_11631_),
    .X(_11632_));
 sky130_fd_sc_hd__inv_4 _28310_ (.A(_11632_),
    .Y(_11633_));
 sky130_fd_sc_hd__a2bb2oi_4 _28311_ (.A1_N(_14286_),
    .A2_N(_11548_),
    .B1(_11547_),
    .B2(_11549_),
    .Y(_11634_));
 sky130_fd_sc_hd__and2_2 _28312_ (.A(_09388_),
    .B(_08492_),
    .X(_11635_));
 sky130_fd_sc_hd__nand3_4 _28313_ (.A(_11132_),
    .B(_10516_),
    .C(_08488_),
    .Y(_11636_));
 sky130_fd_sc_hd__a22o_2 _28314_ (.A1(_07247_),
    .A2(_08073_),
    .B1(_10516_),
    .B2(_08806_),
    .X(_11637_));
 sky130_fd_sc_hd__o21ai_4 _28315_ (.A1(_14280_),
    .A2(_11636_),
    .B1(_11637_),
    .Y(_11638_));
 sky130_fd_sc_hd__xor2_4 _28316_ (.A(_11635_),
    .B(_11638_),
    .X(_11639_));
 sky130_fd_sc_hd__xnor2_4 _28317_ (.A(_11634_),
    .B(_11639_),
    .Y(_11640_));
 sky130_fd_sc_hd__xor2_4 _28318_ (.A(_11633_),
    .B(_11640_),
    .X(_11641_));
 sky130_fd_sc_hd__nor2_1 _28319_ (.A(_11562_),
    .B(_11567_),
    .Y(_11642_));
 sky130_fd_sc_hd__o21bai_2 _28320_ (.A1(_11561_),
    .A2(_11568_),
    .B1_N(_11642_),
    .Y(_11643_));
 sky130_fd_sc_hd__xnor2_2 _28321_ (.A(_11641_),
    .B(_11643_),
    .Y(_11644_));
 sky130_fd_sc_hd__xor2_1 _28322_ (.A(_11629_),
    .B(_11644_),
    .X(_11645_));
 sky130_vsdinv _28323_ (.A(_11645_),
    .Y(_11646_));
 sky130_fd_sc_hd__and2_1 _28324_ (.A(_11585_),
    .B(_11571_),
    .X(_11647_));
 sky130_fd_sc_hd__o21bai_2 _28325_ (.A1(_11569_),
    .A2(_11586_),
    .B1_N(_11647_),
    .Y(_11648_));
 sky130_fd_sc_hd__o21a_2 _28326_ (.A1(_11563_),
    .A2(_11566_),
    .B1(_11564_),
    .X(_11649_));
 sky130_fd_sc_hd__a2bb2oi_4 _28327_ (.A1_N(_14322_),
    .A2_N(_11573_),
    .B1(_11572_),
    .B2(_11574_),
    .Y(_11650_));
 sky130_fd_sc_hd__and2_2 _28328_ (.A(_07107_),
    .B(_10825_),
    .X(_11651_));
 sky130_fd_sc_hd__nand3_4 _28329_ (.A(_11008_),
    .B(_11009_),
    .C(_10827_),
    .Y(_11652_));
 sky130_fd_sc_hd__a22o_2 _28330_ (.A1(_10672_),
    .A2(_07775_),
    .B1(_07103_),
    .B2(_08070_),
    .X(_11653_));
 sky130_fd_sc_hd__o21ai_4 _28331_ (.A1(_14298_),
    .A2(_11652_),
    .B1(_11653_),
    .Y(_11654_));
 sky130_fd_sc_hd__xor2_4 _28332_ (.A(_11651_),
    .B(_11654_),
    .X(_11655_));
 sky130_fd_sc_hd__xnor2_4 _28333_ (.A(_11650_),
    .B(_11655_),
    .Y(_11656_));
 sky130_fd_sc_hd__xnor2_4 _28334_ (.A(_11649_),
    .B(_11656_),
    .Y(_11657_));
 sky130_fd_sc_hd__or2b_1 _28335_ (.A(_11583_),
    .B_N(_11578_),
    .X(_11658_));
 sky130_fd_sc_hd__o21ai_4 _28336_ (.A1(_11576_),
    .A2(_11584_),
    .B1(_11658_),
    .Y(_11659_));
 sky130_fd_sc_hd__and2_2 _28337_ (.A(_07359_),
    .B(_07468_),
    .X(_11660_));
 sky130_fd_sc_hd__nand3_4 _28338_ (.A(_08397_),
    .B(_11020_),
    .C(_08330_),
    .Y(_11661_));
 sky130_fd_sc_hd__a22o_2 _28339_ (.A1(_13972_),
    .A2(_08330_),
    .B1(_11020_),
    .B2(_07473_),
    .X(_11662_));
 sky130_fd_sc_hd__o21ai_4 _28340_ (.A1(_08464_),
    .A2(_11661_),
    .B1(_11662_),
    .Y(_11663_));
 sky130_fd_sc_hd__xor2_4 _28341_ (.A(_11660_),
    .B(_11663_),
    .X(_11664_));
 sky130_fd_sc_hd__nand3b_2 _28342_ (.A_N(_11580_),
    .B(_08527_),
    .C(_14347_),
    .Y(_11665_));
 sky130_fd_sc_hd__o31ai_4 _28343_ (.A1(_11024_),
    .A2(_14334_),
    .A3(_11582_),
    .B1(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__and2_2 _28344_ (.A(_07945_),
    .B(_08701_),
    .X(_11667_));
 sky130_fd_sc_hd__nand2_2 _28345_ (.A(_13961_),
    .B(_06760_),
    .Y(_11668_));
 sky130_fd_sc_hd__and2b_1 _28346_ (.A_N(_07046_),
    .B(_12804_),
    .X(_11669_));
 sky130_fd_sc_hd__xor2_4 _28347_ (.A(_11668_),
    .B(_11669_),
    .X(_11670_));
 sky130_fd_sc_hd__xor2_4 _28348_ (.A(_11667_),
    .B(_11670_),
    .X(_11671_));
 sky130_fd_sc_hd__xor2_4 _28349_ (.A(_11666_),
    .B(_11671_),
    .X(_11672_));
 sky130_fd_sc_hd__xor2_4 _28350_ (.A(_11664_),
    .B(_11672_),
    .X(_11673_));
 sky130_fd_sc_hd__xnor2_4 _28351_ (.A(_11659_),
    .B(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__xor2_4 _28352_ (.A(_11657_),
    .B(_11674_),
    .X(_11675_));
 sky130_fd_sc_hd__xnor2_1 _28353_ (.A(_11648_),
    .B(_11675_),
    .Y(_11676_));
 sky130_fd_sc_hd__xor2_1 _28354_ (.A(_11646_),
    .B(_11676_),
    .X(_11677_));
 sky130_fd_sc_hd__and2_1 _28355_ (.A(_11587_),
    .B(_11560_),
    .X(_11678_));
 sky130_fd_sc_hd__o21ba_1 _28356_ (.A1(_11558_),
    .A2(_11588_),
    .B1_N(_11678_),
    .X(_11679_));
 sky130_fd_sc_hd__or2b_2 _28357_ (.A(_11677_),
    .B_N(_11679_),
    .X(_11680_));
 sky130_fd_sc_hd__or2b_2 _28358_ (.A(_11679_),
    .B_N(_11677_),
    .X(_11681_));
 sky130_fd_sc_hd__and2_1 _28359_ (.A(_11532_),
    .B(_11528_),
    .X(_11682_));
 sky130_fd_sc_hd__o21bai_2 _28360_ (.A1(_11187_),
    .A2(_11533_),
    .B1_N(_11682_),
    .Y(_11683_));
 sky130_fd_sc_hd__o22a_2 _28361_ (.A1(_14033_),
    .A2(_11337_),
    .B1(_11057_),
    .B2(_11336_),
    .X(_11684_));
 sky130_fd_sc_hd__nand3b_1 _28362_ (.A_N(_11543_),
    .B(_10984_),
    .C(_08589_),
    .Y(_11685_));
 sky130_fd_sc_hd__o21a_2 _28363_ (.A1(_11529_),
    .A2(_11544_),
    .B1(_11685_),
    .X(_11686_));
 sky130_fd_sc_hd__xor2_4 _28364_ (.A(_11684_),
    .B(_11686_),
    .X(_11687_));
 sky130_fd_sc_hd__and2_1 _28365_ (.A(_11530_),
    .B(_11339_),
    .X(_11688_));
 sky130_fd_sc_hd__o21bai_4 _28366_ (.A1(_11401_),
    .A2(_11531_),
    .B1_N(_11688_),
    .Y(_11689_));
 sky130_fd_sc_hd__xor2_4 _28367_ (.A(_11687_),
    .B(_11689_),
    .X(_11690_));
 sky130_fd_sc_hd__xor2_4 _28368_ (.A(_11050_),
    .B(_11690_),
    .X(_11691_));
 sky130_fd_sc_hd__and2_1 _28369_ (.A(_11555_),
    .B(_11553_),
    .X(_11692_));
 sky130_fd_sc_hd__o21bai_2 _28370_ (.A1(_11541_),
    .A2(_11556_),
    .B1_N(_11692_),
    .Y(_11693_));
 sky130_fd_sc_hd__xor2_2 _28371_ (.A(_11691_),
    .B(_11693_),
    .X(_11694_));
 sky130_fd_sc_hd__xnor2_2 _28372_ (.A(_11683_),
    .B(_11694_),
    .Y(_11695_));
 sky130_fd_sc_hd__a21oi_1 _28373_ (.A1(_11680_),
    .A2(_11681_),
    .B1(_11695_),
    .Y(_11696_));
 sky130_vsdinv _28374_ (.A(_11696_),
    .Y(_11697_));
 sky130_fd_sc_hd__nand3_4 _28375_ (.A(_11680_),
    .B(_11681_),
    .C(_11695_),
    .Y(_11698_));
 sky130_fd_sc_hd__and2b_1 _28376_ (.A_N(_11539_),
    .B(_11589_),
    .X(_11699_));
 sky130_fd_sc_hd__o21bai_2 _28377_ (.A1(_11537_),
    .A2(_11590_),
    .B1_N(_11699_),
    .Y(_11700_));
 sky130_fd_sc_hd__a21oi_2 _28378_ (.A1(_11697_),
    .A2(_11698_),
    .B1(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__o211a_1 _28379_ (.A1(_11699_),
    .A2(_11591_),
    .B1(_11698_),
    .C1(_11697_),
    .X(_11702_));
 sky130_fd_sc_hd__nand2_1 _28380_ (.A(_11535_),
    .B(_11524_),
    .Y(_11703_));
 sky130_fd_sc_hd__or2_1 _28381_ (.A(_11526_),
    .B(_11534_),
    .X(_11704_));
 sky130_fd_sc_hd__a21o_1 _28382_ (.A1(_11703_),
    .A2(_11704_),
    .B1(_11363_),
    .X(_11705_));
 sky130_fd_sc_hd__nand3_2 _28383_ (.A(_11703_),
    .B(_11476_),
    .C(_11704_),
    .Y(_11706_));
 sky130_fd_sc_hd__nand2_4 _28384_ (.A(_11705_),
    .B(_11706_),
    .Y(_11707_));
 sky130_fd_sc_hd__xor2_4 _28385_ (.A(_11472_),
    .B(_11707_),
    .X(_11708_));
 sky130_fd_sc_hd__o21bai_2 _28386_ (.A1(_11701_),
    .A2(_11702_),
    .B1_N(_11708_),
    .Y(_11709_));
 sky130_fd_sc_hd__nand3b_4 _28387_ (.A_N(_11696_),
    .B(_11700_),
    .C(_11698_),
    .Y(_11710_));
 sky130_fd_sc_hd__nand3b_4 _28388_ (.A_N(_11701_),
    .B(_11710_),
    .C(_11708_),
    .Y(_11711_));
 sky130_fd_sc_hd__o21bai_2 _28389_ (.A1(_11518_),
    .A2(_11594_),
    .B1_N(_11593_),
    .Y(_11712_));
 sky130_fd_sc_hd__a21oi_4 _28390_ (.A1(_11709_),
    .A2(_11711_),
    .B1(_11712_),
    .Y(_11713_));
 sky130_fd_sc_hd__and3_1 _28391_ (.A(_11709_),
    .B(_11711_),
    .C(_11712_),
    .X(_11714_));
 sky130_vsdinv _28392_ (.A(_11714_),
    .Y(_11715_));
 sky130_fd_sc_hd__a21boi_4 _28393_ (.A1(_11602_),
    .A2(_11515_),
    .B1_N(_11514_),
    .Y(_11716_));
 sky130_fd_sc_hd__xor2_4 _28394_ (.A(_10337_),
    .B(_11716_),
    .X(_11717_));
 sky130_fd_sc_hd__nand3b_4 _28395_ (.A_N(_11713_),
    .B(_11715_),
    .C(_11717_),
    .Y(_11718_));
 sky130_fd_sc_hd__o21bai_2 _28396_ (.A1(_11713_),
    .A2(_11714_),
    .B1_N(_11717_),
    .Y(_11719_));
 sky130_vsdinv _28397_ (.A(_11605_),
    .Y(_11720_));
 sky130_fd_sc_hd__a21oi_1 _28398_ (.A1(_11596_),
    .A2(_11597_),
    .B1(_11598_),
    .Y(_11721_));
 sky130_fd_sc_hd__o21ai_2 _28399_ (.A1(_11720_),
    .A2(_11721_),
    .B1(_11600_),
    .Y(_11722_));
 sky130_fd_sc_hd__nand3_4 _28400_ (.A(_11718_),
    .B(_11719_),
    .C(_11722_),
    .Y(_11723_));
 sky130_fd_sc_hd__a21o_1 _28401_ (.A1(_11718_),
    .A2(_11719_),
    .B1(_11722_),
    .X(_11724_));
 sky130_fd_sc_hd__o2bb2ai_1 _28402_ (.A1_N(_11723_),
    .A2_N(_11724_),
    .B1(_11243_),
    .B2(_11604_),
    .Y(_11725_));
 sky130_fd_sc_hd__nor2_1 _28403_ (.A(_10813_),
    .B(_11604_),
    .Y(_11726_));
 sky130_fd_sc_hd__nand3_2 _28404_ (.A(_11724_),
    .B(_11726_),
    .C(_11723_),
    .Y(_11727_));
 sky130_vsdinv _28405_ (.A(_11617_),
    .Y(_11728_));
 sky130_fd_sc_hd__a21oi_1 _28406_ (.A1(_11606_),
    .A2(_11610_),
    .B1(_11609_),
    .Y(_11729_));
 sky130_fd_sc_hd__o21ai_2 _28407_ (.A1(_11728_),
    .A2(_11729_),
    .B1(_11611_),
    .Y(_11730_));
 sky130_fd_sc_hd__a21o_1 _28408_ (.A1(_11725_),
    .A2(_11727_),
    .B1(_11730_),
    .X(_11731_));
 sky130_fd_sc_hd__nand3_2 _28409_ (.A(_11725_),
    .B(_11730_),
    .C(_11727_),
    .Y(_11732_));
 sky130_fd_sc_hd__nand2_1 _28410_ (.A(_11731_),
    .B(_11732_),
    .Y(_11733_));
 sky130_fd_sc_hd__nand3_1 _28411_ (.A(_11620_),
    .B(_11616_),
    .C(_11618_),
    .Y(_11734_));
 sky130_fd_sc_hd__o21ai_2 _28412_ (.A1(_11505_),
    .A2(_11621_),
    .B1(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__a31oi_4 _28413_ (.A1(_11507_),
    .A2(_11626_),
    .A3(_11510_),
    .B1(_11735_),
    .Y(_11736_));
 sky130_vsdinv _28414_ (.A(_11736_),
    .Y(_11737_));
 sky130_fd_sc_hd__a41oi_4 _28415_ (.A1(_11269_),
    .A2(_11507_),
    .A3(_11508_),
    .A4(_11626_),
    .B1(_11737_),
    .Y(_11738_));
 sky130_fd_sc_hd__xor2_1 _28416_ (.A(_11733_),
    .B(_11738_),
    .X(_02671_));
 sky130_fd_sc_hd__or2_1 _28417_ (.A(_11634_),
    .B(_11639_),
    .X(_11739_));
 sky130_fd_sc_hd__o21a_2 _28418_ (.A1(_11633_),
    .A2(_11640_),
    .B1(_11739_),
    .X(_11740_));
 sky130_fd_sc_hd__nor2_1 _28419_ (.A(_11650_),
    .B(_11655_),
    .Y(_11741_));
 sky130_fd_sc_hd__o21bai_4 _28420_ (.A1(_11649_),
    .A2(_11656_),
    .B1_N(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__a2bb2oi_4 _28421_ (.A1_N(_14281_),
    .A2_N(_11636_),
    .B1(_11635_),
    .B2(_11637_),
    .Y(_11743_));
 sky130_fd_sc_hd__nand2_8 _28422_ (.A(_12779_),
    .B(_09388_),
    .Y(_11744_));
 sky130_fd_sc_hd__or4_4 _28423_ (.A(_13999_),
    .B(_14002_),
    .C(_14275_),
    .D(_14279_),
    .X(_11745_));
 sky130_fd_sc_hd__a22o_1 _28424_ (.A1(_11132_),
    .A2(_08480_),
    .B1(_11133_),
    .B2(_08595_),
    .X(_11746_));
 sky130_fd_sc_hd__nand2_4 _28425_ (.A(_11745_),
    .B(_11746_),
    .Y(_11747_));
 sky130_fd_sc_hd__xnor2_4 _28426_ (.A(_11744_),
    .B(_11747_),
    .Y(_11748_));
 sky130_fd_sc_hd__xnor2_4 _28427_ (.A(_11743_),
    .B(_11748_),
    .Y(_11749_));
 sky130_fd_sc_hd__xor2_4 _28428_ (.A(_11633_),
    .B(_11749_),
    .X(_11750_));
 sky130_fd_sc_hd__xnor2_4 _28429_ (.A(_11742_),
    .B(_11750_),
    .Y(_11751_));
 sky130_fd_sc_hd__xor2_2 _28430_ (.A(_11740_),
    .B(_11751_),
    .X(_11752_));
 sky130_fd_sc_hd__and2_1 _28431_ (.A(_11673_),
    .B(_11659_),
    .X(_11753_));
 sky130_fd_sc_hd__o21bai_2 _28432_ (.A1(_11657_),
    .A2(_11674_),
    .B1_N(_11753_),
    .Y(_11754_));
 sky130_fd_sc_hd__a2bb2oi_4 _28433_ (.A1_N(_14300_),
    .A2_N(_11652_),
    .B1(_11651_),
    .B2(_11653_),
    .Y(_11755_));
 sky130_fd_sc_hd__a2bb2oi_4 _28434_ (.A1_N(_14316_),
    .A2_N(_11661_),
    .B1(_11660_),
    .B2(_11662_),
    .Y(_11756_));
 sky130_fd_sc_hd__and2_2 _28435_ (.A(_07107_),
    .B(_08157_),
    .X(_11757_));
 sky130_fd_sc_hd__nand3_4 _28436_ (.A(_11008_),
    .B(_11009_),
    .C(_07769_),
    .Y(_11758_));
 sky130_fd_sc_hd__a22o_2 _28437_ (.A1(_10672_),
    .A2(_08070_),
    .B1(_07103_),
    .B2(_08064_),
    .X(_11759_));
 sky130_fd_sc_hd__o21ai_4 _28438_ (.A1(_14292_),
    .A2(_11758_),
    .B1(_11759_),
    .Y(_11760_));
 sky130_fd_sc_hd__xor2_4 _28439_ (.A(_11757_),
    .B(_11760_),
    .X(_11761_));
 sky130_fd_sc_hd__xnor2_4 _28440_ (.A(_11756_),
    .B(_11761_),
    .Y(_11762_));
 sky130_fd_sc_hd__xnor2_4 _28441_ (.A(_11755_),
    .B(_11762_),
    .Y(_11763_));
 sky130_fd_sc_hd__or2b_1 _28442_ (.A(_11671_),
    .B_N(_11666_),
    .X(_11764_));
 sky130_fd_sc_hd__o21ai_4 _28443_ (.A1(_11664_),
    .A2(_11672_),
    .B1(_11764_),
    .Y(_11765_));
 sky130_fd_sc_hd__and2_2 _28444_ (.A(_07359_),
    .B(_07570_),
    .X(_11766_));
 sky130_fd_sc_hd__nand3_4 _28445_ (.A(_11018_),
    .B(_13979_),
    .C(_07199_),
    .Y(_11767_));
 sky130_fd_sc_hd__a22o_2 _28446_ (.A1(_13972_),
    .A2(_07473_),
    .B1(_11020_),
    .B2(_08885_),
    .X(_11768_));
 sky130_fd_sc_hd__o21ai_4 _28447_ (.A1(_14309_),
    .A2(_11767_),
    .B1(_11768_),
    .Y(_11769_));
 sky130_fd_sc_hd__xor2_4 _28448_ (.A(_11766_),
    .B(_11769_),
    .X(_11770_));
 sky130_fd_sc_hd__nand3b_2 _28449_ (.A_N(_11668_),
    .B(_08527_),
    .C(_14340_),
    .Y(_11771_));
 sky130_fd_sc_hd__o31ai_4 _28450_ (.A1(_11024_),
    .A2(_08332_),
    .A3(_11670_),
    .B1(_11771_),
    .Y(_11772_));
 sky130_fd_sc_hd__and2_2 _28451_ (.A(_11028_),
    .B(_07206_),
    .X(_11773_));
 sky130_fd_sc_hd__nand2_2 _28452_ (.A(_11030_),
    .B(_06596_),
    .Y(_11774_));
 sky130_fd_sc_hd__and2b_1 _28453_ (.A_N(_06760_),
    .B(_12804_),
    .X(_11775_));
 sky130_fd_sc_hd__xor2_4 _28454_ (.A(_11774_),
    .B(_11775_),
    .X(_11776_));
 sky130_fd_sc_hd__xor2_4 _28455_ (.A(_11773_),
    .B(_11776_),
    .X(_11777_));
 sky130_fd_sc_hd__xor2_4 _28456_ (.A(_11772_),
    .B(_11777_),
    .X(_11778_));
 sky130_fd_sc_hd__xor2_4 _28457_ (.A(_11770_),
    .B(_11778_),
    .X(_11779_));
 sky130_fd_sc_hd__xnor2_4 _28458_ (.A(_11765_),
    .B(_11779_),
    .Y(_11780_));
 sky130_fd_sc_hd__xor2_4 _28459_ (.A(_11763_),
    .B(_11780_),
    .X(_11781_));
 sky130_fd_sc_hd__xnor2_1 _28460_ (.A(_11754_),
    .B(_11781_),
    .Y(_11782_));
 sky130_fd_sc_hd__xnor2_1 _28461_ (.A(_11752_),
    .B(_11782_),
    .Y(_11783_));
 sky130_fd_sc_hd__and2_1 _28462_ (.A(_11675_),
    .B(_11648_),
    .X(_11784_));
 sky130_fd_sc_hd__o21ba_1 _28463_ (.A1(_11646_),
    .A2(_11676_),
    .B1_N(_11784_),
    .X(_11785_));
 sky130_fd_sc_hd__or2b_2 _28464_ (.A(_11783_),
    .B_N(_11785_),
    .X(_11786_));
 sky130_fd_sc_hd__or2b_4 _28465_ (.A(_11785_),
    .B_N(_11783_),
    .X(_11787_));
 sky130_fd_sc_hd__or2b_1 _28466_ (.A(_11687_),
    .B_N(_11689_),
    .X(_11788_));
 sky130_fd_sc_hd__o21a_4 _28467_ (.A1(_11187_),
    .A2(_11690_),
    .B1(_11788_),
    .X(_11789_));
 sky130_fd_sc_hd__o22a_4 _28468_ (.A1(_14011_),
    .A2(_11543_),
    .B1(_11529_),
    .B2(_11631_),
    .X(_11790_));
 sky130_fd_sc_hd__o31a_1 _28469_ (.A1(_07295_),
    .A2(_05815_),
    .A3(_05718_),
    .B1(_12781_),
    .X(_11791_));
 sky130_fd_sc_hd__nand3b_4 _28470_ (.A_N(_11197_),
    .B(_07295_),
    .C(_05718_),
    .Y(_11792_));
 sky130_fd_sc_hd__a21boi_4 _28471_ (.A1(_11686_),
    .A2(_11791_),
    .B1_N(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__xor2_4 _28472_ (.A(_11790_),
    .B(_11793_),
    .X(_11794_));
 sky130_fd_sc_hd__xnor2_4 _28473_ (.A(_11050_),
    .B(_11794_),
    .Y(_11795_));
 sky130_fd_sc_hd__and2_1 _28474_ (.A(_11643_),
    .B(_11641_),
    .X(_11796_));
 sky130_fd_sc_hd__o21bai_4 _28475_ (.A1(_11629_),
    .A2(_11644_),
    .B1_N(_11796_),
    .Y(_11797_));
 sky130_fd_sc_hd__xor2_4 _28476_ (.A(_11795_),
    .B(_11797_),
    .X(_11798_));
 sky130_fd_sc_hd__xor2_4 _28477_ (.A(_11789_),
    .B(_11798_),
    .X(_11799_));
 sky130_fd_sc_hd__a21o_1 _28478_ (.A1(_11786_),
    .A2(_11787_),
    .B1(_11799_),
    .X(_11800_));
 sky130_fd_sc_hd__nand3_4 _28479_ (.A(_11786_),
    .B(_11787_),
    .C(_11799_),
    .Y(_11801_));
 sky130_fd_sc_hd__nand2_2 _28480_ (.A(_11698_),
    .B(_11681_),
    .Y(_11802_));
 sky130_fd_sc_hd__a21oi_4 _28481_ (.A1(_11800_),
    .A2(_11801_),
    .B1(_11802_),
    .Y(_11803_));
 sky130_vsdinv _28482_ (.A(_11803_),
    .Y(_11804_));
 sky130_fd_sc_hd__nand3_4 _28483_ (.A(_11802_),
    .B(_11800_),
    .C(_11801_),
    .Y(_11805_));
 sky130_fd_sc_hd__and2b_1 _28484_ (.A_N(_11691_),
    .B(_11693_),
    .X(_11806_));
 sky130_fd_sc_hd__and2b_1 _28485_ (.A_N(_11694_),
    .B(_11683_),
    .X(_11807_));
 sky130_fd_sc_hd__or3_4 _28486_ (.A(_11361_),
    .B(_11806_),
    .C(_11807_),
    .X(_11808_));
 sky130_fd_sc_hd__o21bai_1 _28487_ (.A1(_11806_),
    .A2(_11807_),
    .B1_N(_11363_),
    .Y(_11809_));
 sky130_fd_sc_hd__nand2_2 _28488_ (.A(_11808_),
    .B(_11809_),
    .Y(_11810_));
 sky130_fd_sc_hd__xor2_4 _28489_ (.A(_11601_),
    .B(_11810_),
    .X(_11811_));
 sky130_fd_sc_hd__a21bo_1 _28490_ (.A1(_11804_),
    .A2(_11805_),
    .B1_N(_11811_),
    .X(_11812_));
 sky130_fd_sc_hd__nand3b_4 _28491_ (.A_N(_11811_),
    .B(_11804_),
    .C(_11805_),
    .Y(_11813_));
 sky130_fd_sc_hd__nand2_2 _28492_ (.A(_11711_),
    .B(_11710_),
    .Y(_11814_));
 sky130_fd_sc_hd__a21o_1 _28493_ (.A1(_11812_),
    .A2(_11813_),
    .B1(_11814_),
    .X(_11815_));
 sky130_fd_sc_hd__nand3_4 _28494_ (.A(_11814_),
    .B(_11813_),
    .C(_11812_),
    .Y(_11816_));
 sky130_fd_sc_hd__o21ai_4 _28495_ (.A1(_11473_),
    .A2(_11707_),
    .B1(_11705_),
    .Y(_11817_));
 sky130_fd_sc_hd__xor2_4 _28496_ (.A(_10178_),
    .B(_11817_),
    .X(_11818_));
 sky130_fd_sc_hd__a21oi_2 _28497_ (.A1(_11815_),
    .A2(_11816_),
    .B1(_11818_),
    .Y(_11819_));
 sky130_fd_sc_hd__nand3_4 _28498_ (.A(_11815_),
    .B(_11816_),
    .C(_11818_),
    .Y(_11820_));
 sky130_vsdinv _28499_ (.A(_11717_),
    .Y(_11821_));
 sky130_fd_sc_hd__o21bai_2 _28500_ (.A1(_11713_),
    .A2(_11821_),
    .B1_N(_11714_),
    .Y(_11822_));
 sky130_fd_sc_hd__nand3b_4 _28501_ (.A_N(_11819_),
    .B(_11820_),
    .C(_11822_),
    .Y(_11823_));
 sky130_vsdinv _28502_ (.A(_11820_),
    .Y(_11824_));
 sky130_fd_sc_hd__o21bai_2 _28503_ (.A1(_11819_),
    .A2(_11824_),
    .B1_N(_11822_),
    .Y(_11825_));
 sky130_fd_sc_hd__o2bb2ai_1 _28504_ (.A1_N(_11823_),
    .A2_N(_11825_),
    .B1(_11243_),
    .B2(_11716_),
    .Y(_11826_));
 sky130_fd_sc_hd__nor2_2 _28505_ (.A(_11242_),
    .B(_11716_),
    .Y(_11827_));
 sky130_fd_sc_hd__nand3_4 _28506_ (.A(_11825_),
    .B(_11823_),
    .C(_11827_),
    .Y(_11828_));
 sky130_vsdinv _28507_ (.A(_11726_),
    .Y(_11829_));
 sky130_fd_sc_hd__a21oi_1 _28508_ (.A1(_11718_),
    .A2(_11719_),
    .B1(_11722_),
    .Y(_11830_));
 sky130_fd_sc_hd__o21ai_2 _28509_ (.A1(_11829_),
    .A2(_11830_),
    .B1(_11723_),
    .Y(_11831_));
 sky130_fd_sc_hd__a21o_1 _28510_ (.A1(_11826_),
    .A2(_11828_),
    .B1(_11831_),
    .X(_11832_));
 sky130_fd_sc_hd__nand3_1 _28511_ (.A(_11826_),
    .B(_11831_),
    .C(_11828_),
    .Y(_11833_));
 sky130_fd_sc_hd__nand2_1 _28512_ (.A(_11832_),
    .B(_11833_),
    .Y(_11834_));
 sky130_fd_sc_hd__o21ai_1 _28513_ (.A1(_11733_),
    .A2(_11738_),
    .B1(_11732_),
    .Y(_11835_));
 sky130_fd_sc_hd__xnor2_1 _28514_ (.A(_11834_),
    .B(_11835_),
    .Y(_02672_));
 sky130_fd_sc_hd__or2_1 _28515_ (.A(_11743_),
    .B(_11748_),
    .X(_11836_));
 sky130_fd_sc_hd__o21a_1 _28516_ (.A1(_11633_),
    .A2(_11749_),
    .B1(_11836_),
    .X(_11837_));
 sky130_fd_sc_hd__or2_1 _28517_ (.A(_11756_),
    .B(_11761_),
    .X(_11838_));
 sky130_fd_sc_hd__o21a_1 _28518_ (.A1(_11755_),
    .A2(_11762_),
    .B1(_11838_),
    .X(_11839_));
 sky130_fd_sc_hd__clkbuf_8 _28519_ (.A(_11632_),
    .X(_11840_));
 sky130_fd_sc_hd__nand3_4 _28520_ (.A(_12779_),
    .B(_11132_),
    .C(_08595_),
    .Y(_11841_));
 sky130_fd_sc_hd__a22o_2 _28521_ (.A1(_09283_),
    .A2(_10516_),
    .B1(_10515_),
    .B2(_08595_),
    .X(_11842_));
 sky130_fd_sc_hd__o21ai_4 _28522_ (.A1(_14002_),
    .A2(_11841_),
    .B1(_11842_),
    .Y(_11843_));
 sky130_fd_sc_hd__xor2_4 _28523_ (.A(_11744_),
    .B(_11843_),
    .X(_11844_));
 sky130_fd_sc_hd__o21ai_4 _28524_ (.A1(_11744_),
    .A2(_11747_),
    .B1(_11745_),
    .Y(_11845_));
 sky130_fd_sc_hd__xnor2_4 _28525_ (.A(_11844_),
    .B(_11845_),
    .Y(_11846_));
 sky130_fd_sc_hd__xor2_4 _28526_ (.A(_11840_),
    .B(_11846_),
    .X(_11847_));
 sky130_fd_sc_hd__xnor2_2 _28527_ (.A(_11839_),
    .B(_11847_),
    .Y(_11848_));
 sky130_fd_sc_hd__xor2_1 _28528_ (.A(_11837_),
    .B(_11848_),
    .X(_11849_));
 sky130_vsdinv _28529_ (.A(_11849_),
    .Y(_11850_));
 sky130_fd_sc_hd__and2_1 _28530_ (.A(_11779_),
    .B(_11765_),
    .X(_11851_));
 sky130_fd_sc_hd__o21bai_2 _28531_ (.A1(_11763_),
    .A2(_11780_),
    .B1_N(_11851_),
    .Y(_11852_));
 sky130_fd_sc_hd__a2bb2oi_4 _28532_ (.A1_N(_14294_),
    .A2_N(_11758_),
    .B1(_11757_),
    .B2(_11759_),
    .Y(_11853_));
 sky130_fd_sc_hd__a2bb2oi_4 _28533_ (.A1_N(_14311_),
    .A2_N(_11767_),
    .B1(_11766_),
    .B2(_11768_),
    .Y(_11854_));
 sky130_fd_sc_hd__nand2_2 _28534_ (.A(net437),
    .B(_08481_),
    .Y(_11855_));
 sky130_fd_sc_hd__or4_4 _28535_ (.A(_13986_),
    .B(_13991_),
    .C(_08084_),
    .D(_14291_),
    .X(_11856_));
 sky130_fd_sc_hd__a22o_1 _28536_ (.A1(_11008_),
    .A2(_08064_),
    .B1(_11009_),
    .B2(_08157_),
    .X(_11857_));
 sky130_fd_sc_hd__nand2_2 _28537_ (.A(_11856_),
    .B(_11857_),
    .Y(_11858_));
 sky130_fd_sc_hd__xnor2_4 _28538_ (.A(_11855_),
    .B(_11858_),
    .Y(_11859_));
 sky130_fd_sc_hd__xnor2_4 _28539_ (.A(_11854_),
    .B(_11859_),
    .Y(_11860_));
 sky130_fd_sc_hd__xnor2_4 _28540_ (.A(_11853_),
    .B(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__or2b_2 _28541_ (.A(_11777_),
    .B_N(_11772_),
    .X(_11862_));
 sky130_fd_sc_hd__o21ai_4 _28542_ (.A1(_11770_),
    .A2(_11778_),
    .B1(_11862_),
    .Y(_11863_));
 sky130_fd_sc_hd__and2_2 _28543_ (.A(_11162_),
    .B(_10829_),
    .X(_11864_));
 sky130_fd_sc_hd__nand3_4 _28544_ (.A(_11018_),
    .B(_11166_),
    .C(_07468_),
    .Y(_11865_));
 sky130_fd_sc_hd__a22o_2 _28545_ (.A1(_08397_),
    .A2(_07575_),
    .B1(_13979_),
    .B2(_10827_),
    .X(_11866_));
 sky130_fd_sc_hd__o21ai_4 _28546_ (.A1(_09222_),
    .A2(_11865_),
    .B1(_11866_),
    .Y(_11867_));
 sky130_fd_sc_hd__xor2_4 _28547_ (.A(_11864_),
    .B(_11867_),
    .X(_11868_));
 sky130_fd_sc_hd__nand3b_4 _28548_ (.A_N(_11774_),
    .B(_11025_),
    .C(_14334_),
    .Y(_11869_));
 sky130_fd_sc_hd__o31ai_4 _28549_ (.A1(_11024_),
    .A2(_14321_),
    .A3(_11776_),
    .B1(_11869_),
    .Y(_11870_));
 sky130_fd_sc_hd__and2_2 _28550_ (.A(_11028_),
    .B(_07198_),
    .X(_11871_));
 sky130_fd_sc_hd__nand2_2 _28551_ (.A(_11030_),
    .B(_07205_),
    .Y(_11872_));
 sky130_fd_sc_hd__and2b_2 _28552_ (.A_N(_06596_),
    .B(_12805_),
    .X(_11873_));
 sky130_fd_sc_hd__xor2_4 _28553_ (.A(_11872_),
    .B(_11873_),
    .X(_11874_));
 sky130_fd_sc_hd__xor2_4 _28554_ (.A(_11871_),
    .B(_11874_),
    .X(_11875_));
 sky130_fd_sc_hd__xor2_4 _28555_ (.A(_11870_),
    .B(_11875_),
    .X(_11876_));
 sky130_fd_sc_hd__xor2_4 _28556_ (.A(_11868_),
    .B(_11876_),
    .X(_11877_));
 sky130_fd_sc_hd__xnor2_4 _28557_ (.A(_11863_),
    .B(_11877_),
    .Y(_11878_));
 sky130_fd_sc_hd__xor2_2 _28558_ (.A(_11861_),
    .B(_11878_),
    .X(_11879_));
 sky130_fd_sc_hd__xnor2_1 _28559_ (.A(_11852_),
    .B(_11879_),
    .Y(_11880_));
 sky130_fd_sc_hd__xor2_1 _28560_ (.A(_11850_),
    .B(_11880_),
    .X(_11881_));
 sky130_fd_sc_hd__or2_1 _28561_ (.A(_11754_),
    .B(_11781_),
    .X(_11882_));
 sky130_fd_sc_hd__and2_1 _28562_ (.A(_11781_),
    .B(_11754_),
    .X(_11883_));
 sky130_fd_sc_hd__a21oi_1 _28563_ (.A1(_11882_),
    .A2(_11752_),
    .B1(_11883_),
    .Y(_11884_));
 sky130_fd_sc_hd__or2b_2 _28564_ (.A(_11881_),
    .B_N(_11884_),
    .X(_11885_));
 sky130_fd_sc_hd__or2b_4 _28565_ (.A(_11884_),
    .B_N(_11881_),
    .X(_11886_));
 sky130_fd_sc_hd__nor2_8 _28566_ (.A(_11792_),
    .B(_11790_),
    .Y(_11887_));
 sky130_fd_sc_hd__a21oi_4 _28567_ (.A1(_11794_),
    .A2(_11330_),
    .B1(_11887_),
    .Y(_11888_));
 sky130_fd_sc_hd__nand3b_4 _28568_ (.A_N(_11336_),
    .B(_11790_),
    .C(_11333_),
    .Y(_11889_));
 sky130_fd_sc_hd__o21ai_4 _28569_ (.A1(_11792_),
    .A2(_11790_),
    .B1(_11889_),
    .Y(_11890_));
 sky130_fd_sc_hd__xnor2_4 _28570_ (.A(_11890_),
    .B(_11050_),
    .Y(_11891_));
 sky130_fd_sc_hd__clkinv_4 _28571_ (.A(_11891_),
    .Y(_11892_));
 sky130_fd_sc_hd__and2_1 _28572_ (.A(_11750_),
    .B(_11742_),
    .X(_11893_));
 sky130_fd_sc_hd__o21bai_4 _28573_ (.A1(_11740_),
    .A2(_11751_),
    .B1_N(_11893_),
    .Y(_11894_));
 sky130_fd_sc_hd__xor2_4 _28574_ (.A(_11892_),
    .B(_11894_),
    .X(_11895_));
 sky130_fd_sc_hd__xor2_4 _28575_ (.A(_11888_),
    .B(_11895_),
    .X(_11896_));
 sky130_fd_sc_hd__a21oi_4 _28576_ (.A1(_11885_),
    .A2(_11886_),
    .B1(_11896_),
    .Y(_11897_));
 sky130_vsdinv _28577_ (.A(_11897_),
    .Y(_11898_));
 sky130_fd_sc_hd__nand3_4 _28578_ (.A(_11885_),
    .B(_11886_),
    .C(_11896_),
    .Y(_11899_));
 sky130_fd_sc_hd__nand2_4 _28579_ (.A(_11801_),
    .B(_11787_),
    .Y(_11900_));
 sky130_fd_sc_hd__a21oi_4 _28580_ (.A1(_11898_),
    .A2(_11899_),
    .B1(_11900_),
    .Y(_11901_));
 sky130_fd_sc_hd__nand3b_4 _28581_ (.A_N(_11897_),
    .B(_11899_),
    .C(_11900_),
    .Y(_11902_));
 sky130_fd_sc_hd__or2_1 _28582_ (.A(_11789_),
    .B(_11798_),
    .X(_11903_));
 sky130_fd_sc_hd__or2b_2 _28583_ (.A(_11795_),
    .B_N(_11797_),
    .X(_11904_));
 sky130_fd_sc_hd__a21o_1 _28584_ (.A1(_11903_),
    .A2(_11904_),
    .B1(_11363_),
    .X(_11905_));
 sky130_fd_sc_hd__o211ai_4 _28585_ (.A1(_11789_),
    .A2(_11798_),
    .B1(_11363_),
    .C1(_11904_),
    .Y(_11906_));
 sky130_fd_sc_hd__a21oi_4 _28586_ (.A1(_11905_),
    .A2(_11906_),
    .B1(_11601_),
    .Y(_11907_));
 sky130_fd_sc_hd__o211a_1 _28587_ (.A1(_11353_),
    .A2(_11357_),
    .B1(_11906_),
    .C1(_11905_),
    .X(_11908_));
 sky130_fd_sc_hd__nor2_2 _28588_ (.A(_11907_),
    .B(_11908_),
    .Y(_11909_));
 sky130_fd_sc_hd__nand3b_4 _28589_ (.A_N(_11901_),
    .B(_11902_),
    .C(_11909_),
    .Y(_11910_));
 sky130_vsdinv _28590_ (.A(_11899_),
    .Y(_11911_));
 sky130_fd_sc_hd__nor3b_4 _28591_ (.A(_11897_),
    .B(_11911_),
    .C_N(_11900_),
    .Y(_11912_));
 sky130_fd_sc_hd__o21bai_4 _28592_ (.A1(_11912_),
    .A2(_11901_),
    .B1_N(_11909_),
    .Y(_11913_));
 sky130_fd_sc_hd__o21ai_4 _28593_ (.A1(_11803_),
    .A2(_11811_),
    .B1(_11805_),
    .Y(_11914_));
 sky130_fd_sc_hd__a21oi_4 _28594_ (.A1(_11910_),
    .A2(_11913_),
    .B1(_11914_),
    .Y(_11915_));
 sky130_fd_sc_hd__and3_1 _28595_ (.A(_11910_),
    .B(_11913_),
    .C(_11914_),
    .X(_11916_));
 sky130_fd_sc_hd__a21boi_4 _28596_ (.A1(_11808_),
    .A2(_11602_),
    .B1_N(_11809_),
    .Y(_11917_));
 sky130_fd_sc_hd__xor2_1 _28597_ (.A(_10325_),
    .B(_11917_),
    .X(_11918_));
 sky130_vsdinv _28598_ (.A(_11918_),
    .Y(_11919_));
 sky130_fd_sc_hd__o21a_1 _28599_ (.A1(_11915_),
    .A2(_11916_),
    .B1(_11919_),
    .X(_11920_));
 sky130_fd_sc_hd__nand3_2 _28600_ (.A(_11910_),
    .B(_11913_),
    .C(_11914_),
    .Y(_11921_));
 sky130_fd_sc_hd__nor3b_4 _28601_ (.A(_11919_),
    .B(_11915_),
    .C_N(_11921_),
    .Y(_11922_));
 sky130_vsdinv _28602_ (.A(_11922_),
    .Y(_11923_));
 sky130_vsdinv _28603_ (.A(_11818_),
    .Y(_11924_));
 sky130_fd_sc_hd__a21oi_1 _28604_ (.A1(_11812_),
    .A2(_11813_),
    .B1(_11814_),
    .Y(_11925_));
 sky130_fd_sc_hd__o21ai_2 _28605_ (.A1(_11924_),
    .A2(_11925_),
    .B1(_11816_),
    .Y(_11926_));
 sky130_fd_sc_hd__nand3b_4 _28606_ (.A_N(_11920_),
    .B(_11923_),
    .C(_11926_),
    .Y(_11927_));
 sky130_fd_sc_hd__o21bai_2 _28607_ (.A1(_11922_),
    .A2(_11920_),
    .B1_N(_11926_),
    .Y(_11928_));
 sky130_fd_sc_hd__and2_1 _28608_ (.A(_11817_),
    .B(_10178_),
    .X(_11929_));
 sky130_fd_sc_hd__a21o_1 _28609_ (.A1(_11927_),
    .A2(_11928_),
    .B1(_11929_),
    .X(_11930_));
 sky130_fd_sc_hd__nand3_2 _28610_ (.A(_11927_),
    .B(_11929_),
    .C(_11928_),
    .Y(_11931_));
 sky130_fd_sc_hd__nand2_1 _28611_ (.A(_11828_),
    .B(_11823_),
    .Y(_11932_));
 sky130_fd_sc_hd__a21oi_2 _28612_ (.A1(_11930_),
    .A2(_11931_),
    .B1(_11932_),
    .Y(_11933_));
 sky130_fd_sc_hd__nand2_1 _28613_ (.A(_11930_),
    .B(_11931_),
    .Y(_11934_));
 sky130_fd_sc_hd__a21oi_4 _28614_ (.A1(_11823_),
    .A2(_11828_),
    .B1(_11934_),
    .Y(_11935_));
 sky130_fd_sc_hd__nor2_2 _28615_ (.A(_11933_),
    .B(_11935_),
    .Y(_11936_));
 sky130_fd_sc_hd__nor2_1 _28616_ (.A(_11834_),
    .B(_11733_),
    .Y(_11937_));
 sky130_vsdinv _28617_ (.A(_11937_),
    .Y(_11938_));
 sky130_fd_sc_hd__a21oi_1 _28618_ (.A1(_11826_),
    .A2(_11828_),
    .B1(_11831_),
    .Y(_11939_));
 sky130_fd_sc_hd__a21oi_1 _28619_ (.A1(_11732_),
    .A2(_11833_),
    .B1(_11939_),
    .Y(_11940_));
 sky130_fd_sc_hd__o21bai_1 _28620_ (.A1(_11938_),
    .A2(_11738_),
    .B1_N(_11940_),
    .Y(_11941_));
 sky130_fd_sc_hd__xor2_1 _28621_ (.A(_11936_),
    .B(_11941_),
    .X(_02673_));
 sky130_fd_sc_hd__a21oi_2 _28622_ (.A1(_11330_),
    .A2(_11889_),
    .B1(_11887_),
    .Y(_11942_));
 sky130_vsdinv _28623_ (.A(_11942_),
    .Y(_11943_));
 sky130_fd_sc_hd__nor2_1 _28624_ (.A(_11839_),
    .B(_11847_),
    .Y(_11944_));
 sky130_fd_sc_hd__o21bai_4 _28625_ (.A1(_11837_),
    .A2(_11848_),
    .B1_N(_11944_),
    .Y(_11945_));
 sky130_fd_sc_hd__xor2_4 _28626_ (.A(_11892_),
    .B(_11945_),
    .X(_11946_));
 sky130_fd_sc_hd__xor2_4 _28627_ (.A(_11943_),
    .B(_11946_),
    .X(_11947_));
 sky130_fd_sc_hd__and2_1 _28628_ (.A(_11879_),
    .B(_11852_),
    .X(_11948_));
 sky130_fd_sc_hd__o21ba_2 _28629_ (.A1(_11850_),
    .A2(_11880_),
    .B1_N(_11948_),
    .X(_11949_));
 sky130_fd_sc_hd__nand2_1 _28630_ (.A(_11845_),
    .B(_11844_),
    .Y(_11950_));
 sky130_fd_sc_hd__o21a_2 _28631_ (.A1(_11633_),
    .A2(_11846_),
    .B1(_11950_),
    .X(_11951_));
 sky130_fd_sc_hd__o21ai_2 _28632_ (.A1(_10991_),
    .A2(_10992_),
    .B1(_12780_),
    .Y(_11952_));
 sky130_fd_sc_hd__nand3_4 _28633_ (.A(_12780_),
    .B(_10991_),
    .C(_10992_),
    .Y(_11953_));
 sky130_fd_sc_hd__and2b_2 _28634_ (.A_N(_11952_),
    .B(_11953_),
    .X(_11954_));
 sky130_fd_sc_hd__or2b_1 _28635_ (.A(_11841_),
    .B_N(_10992_),
    .X(_11955_));
 sky130_fd_sc_hd__a22oi_4 _28636_ (.A1(_11842_),
    .A2(_06472_),
    .B1(_11955_),
    .B2(_11744_),
    .Y(_11956_));
 sky130_fd_sc_hd__xor2_4 _28637_ (.A(_11954_),
    .B(_11956_),
    .X(_11957_));
 sky130_fd_sc_hd__xnor2_4 _28638_ (.A(_11840_),
    .B(_11957_),
    .Y(_11958_));
 sky130_fd_sc_hd__or2_1 _28639_ (.A(_11854_),
    .B(_11859_),
    .X(_11959_));
 sky130_fd_sc_hd__o21a_2 _28640_ (.A1(_11853_),
    .A2(_11860_),
    .B1(_11959_),
    .X(_11960_));
 sky130_fd_sc_hd__xnor2_4 _28641_ (.A(_11958_),
    .B(_11960_),
    .Y(_11961_));
 sky130_fd_sc_hd__xor2_4 _28642_ (.A(_11951_),
    .B(_11961_),
    .X(_11962_));
 sky130_fd_sc_hd__and2_1 _28643_ (.A(_11877_),
    .B(_11863_),
    .X(_11963_));
 sky130_fd_sc_hd__o21bai_4 _28644_ (.A1(_11861_),
    .A2(_11878_),
    .B1_N(_11963_),
    .Y(_11964_));
 sky130_fd_sc_hd__o21a_2 _28645_ (.A1(_11855_),
    .A2(_11858_),
    .B1(_11856_),
    .X(_11965_));
 sky130_fd_sc_hd__a2bb2oi_4 _28646_ (.A1_N(_14305_),
    .A2_N(_11865_),
    .B1(_11864_),
    .B2(_11866_),
    .Y(_11966_));
 sky130_fd_sc_hd__nand2_2 _28647_ (.A(net437),
    .B(_08588_),
    .Y(_11967_));
 sky130_fd_sc_hd__or4_4 _28648_ (.A(_13986_),
    .B(_13991_),
    .C(_14280_),
    .D(_08084_),
    .X(_11968_));
 sky130_fd_sc_hd__a22o_1 _28649_ (.A1(_11006_),
    .A2(_08157_),
    .B1(_07104_),
    .B2(_11138_),
    .X(_11969_));
 sky130_fd_sc_hd__nand2_2 _28650_ (.A(_11968_),
    .B(_11969_),
    .Y(_11970_));
 sky130_fd_sc_hd__xnor2_4 _28651_ (.A(_11967_),
    .B(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__xnor2_4 _28652_ (.A(_11966_),
    .B(_11971_),
    .Y(_11972_));
 sky130_fd_sc_hd__xnor2_4 _28653_ (.A(_11965_),
    .B(_11972_),
    .Y(_11973_));
 sky130_fd_sc_hd__or2b_2 _28654_ (.A(_11875_),
    .B_N(_11870_),
    .X(_11974_));
 sky130_fd_sc_hd__o21ai_4 _28655_ (.A1(_11868_),
    .A2(_11876_),
    .B1(_11974_),
    .Y(_11975_));
 sky130_fd_sc_hd__and2_2 _28656_ (.A(_07360_),
    .B(_08065_),
    .X(_11976_));
 sky130_fd_sc_hd__nand3_4 _28657_ (.A(_13973_),
    .B(_11164_),
    .C(_07570_),
    .Y(_11977_));
 sky130_fd_sc_hd__a22o_2 _28658_ (.A1(_13973_),
    .A2(_10827_),
    .B1(_11166_),
    .B2(_10829_),
    .X(_11978_));
 sky130_fd_sc_hd__o21ai_4 _28659_ (.A1(_14299_),
    .A2(_11977_),
    .B1(_11978_),
    .Y(_11979_));
 sky130_fd_sc_hd__xor2_4 _28660_ (.A(_11976_),
    .B(_11979_),
    .X(_11980_));
 sky130_fd_sc_hd__nand3b_2 _28661_ (.A_N(_11872_),
    .B(_08528_),
    .C(_08332_),
    .Y(_11981_));
 sky130_fd_sc_hd__o31ai_4 _28662_ (.A1(_13968_),
    .A2(_08464_),
    .A3(_11874_),
    .B1(_11981_),
    .Y(_11982_));
 sky130_fd_sc_hd__and2_2 _28663_ (.A(_07946_),
    .B(_08885_),
    .X(_11983_));
 sky130_fd_sc_hd__nand2_2 _28664_ (.A(_13962_),
    .B(_07198_),
    .Y(_11984_));
 sky130_fd_sc_hd__and2b_2 _28665_ (.A_N(_07036_),
    .B(_09025_),
    .X(_11985_));
 sky130_fd_sc_hd__xor2_4 _28666_ (.A(_11984_),
    .B(_11985_),
    .X(_11986_));
 sky130_fd_sc_hd__xor2_4 _28667_ (.A(_11983_),
    .B(_11986_),
    .X(_11987_));
 sky130_fd_sc_hd__xor2_4 _28668_ (.A(_11982_),
    .B(_11987_),
    .X(_11988_));
 sky130_fd_sc_hd__xor2_4 _28669_ (.A(_11980_),
    .B(_11988_),
    .X(_11989_));
 sky130_fd_sc_hd__xnor2_4 _28670_ (.A(_11975_),
    .B(_11989_),
    .Y(_11990_));
 sky130_fd_sc_hd__xor2_4 _28671_ (.A(_11973_),
    .B(_11990_),
    .X(_11991_));
 sky130_fd_sc_hd__xnor2_4 _28672_ (.A(_11964_),
    .B(_11991_),
    .Y(_11992_));
 sky130_fd_sc_hd__xnor2_4 _28673_ (.A(_11962_),
    .B(_11992_),
    .Y(_11993_));
 sky130_fd_sc_hd__xor2_4 _28674_ (.A(_11949_),
    .B(_11993_),
    .X(_11994_));
 sky130_fd_sc_hd__nor2_1 _28675_ (.A(_11947_),
    .B(_11994_),
    .Y(_11995_));
 sky130_vsdinv _28676_ (.A(_11995_),
    .Y(_11996_));
 sky130_fd_sc_hd__nand2_2 _28677_ (.A(_11994_),
    .B(_11947_),
    .Y(_11997_));
 sky130_fd_sc_hd__nand2_2 _28678_ (.A(_11899_),
    .B(_11886_),
    .Y(_11998_));
 sky130_fd_sc_hd__a21oi_4 _28679_ (.A1(_11996_),
    .A2(_11997_),
    .B1(_11998_),
    .Y(_11999_));
 sky130_fd_sc_hd__nand3b_4 _28680_ (.A_N(_11995_),
    .B(_11997_),
    .C(_11998_),
    .Y(_12000_));
 sky130_vsdinv _28681_ (.A(_12000_),
    .Y(_12001_));
 sky130_fd_sc_hd__clkbuf_2 _28682_ (.A(_11891_),
    .X(_12002_));
 sky130_fd_sc_hd__nand2_2 _28683_ (.A(_11894_),
    .B(_12002_),
    .Y(_12003_));
 sky130_fd_sc_hd__o211a_2 _28684_ (.A1(_11888_),
    .A2(_11895_),
    .B1(_11476_),
    .C1(_12003_),
    .X(_12004_));
 sky130_fd_sc_hd__or2_1 _28685_ (.A(_11888_),
    .B(_11895_),
    .X(_12005_));
 sky130_fd_sc_hd__a21oi_4 _28686_ (.A1(_12005_),
    .A2(_12003_),
    .B1(_11476_),
    .Y(_12006_));
 sky130_fd_sc_hd__nor3_4 _28687_ (.A(_11473_),
    .B(_12004_),
    .C(_12006_),
    .Y(_12007_));
 sky130_fd_sc_hd__o21a_1 _28688_ (.A1(_12004_),
    .A2(_12006_),
    .B1(_11472_),
    .X(_12008_));
 sky130_fd_sc_hd__nor2_2 _28689_ (.A(_12007_),
    .B(_12008_),
    .Y(_12009_));
 sky130_fd_sc_hd__o21bai_2 _28690_ (.A1(_11999_),
    .A2(_12001_),
    .B1_N(_12009_),
    .Y(_12010_));
 sky130_fd_sc_hd__nand3b_4 _28691_ (.A_N(_11999_),
    .B(_12000_),
    .C(_12009_),
    .Y(_12011_));
 sky130_fd_sc_hd__o31ai_4 _28692_ (.A1(_11908_),
    .A2(_11907_),
    .A3(_11901_),
    .B1(_11902_),
    .Y(_12012_));
 sky130_fd_sc_hd__a21o_1 _28693_ (.A1(_12010_),
    .A2(_12011_),
    .B1(_12012_),
    .X(_12013_));
 sky130_fd_sc_hd__nand3_4 _28694_ (.A(_12012_),
    .B(_12011_),
    .C(_12010_),
    .Y(_12014_));
 sky130_fd_sc_hd__a21boi_4 _28695_ (.A1(_11602_),
    .A2(_11906_),
    .B1_N(_11905_),
    .Y(_12015_));
 sky130_fd_sc_hd__xor2_4 _28696_ (.A(_10337_),
    .B(_12015_),
    .X(_12016_));
 sky130_fd_sc_hd__a21oi_2 _28697_ (.A1(_12013_),
    .A2(_12014_),
    .B1(_12016_),
    .Y(_12017_));
 sky130_fd_sc_hd__nand3_4 _28698_ (.A(_12013_),
    .B(_12014_),
    .C(_12016_),
    .Y(_12018_));
 sky130_fd_sc_hd__o21ai_2 _28699_ (.A1(_11919_),
    .A2(_11915_),
    .B1(_11921_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand3b_4 _28700_ (.A_N(_12017_),
    .B(_12018_),
    .C(_12019_),
    .Y(_12020_));
 sky130_vsdinv _28701_ (.A(_12018_),
    .Y(_12021_));
 sky130_fd_sc_hd__o21bai_2 _28702_ (.A1(_12017_),
    .A2(_12021_),
    .B1_N(_12019_),
    .Y(_12022_));
 sky130_fd_sc_hd__o2bb2ai_1 _28703_ (.A1_N(_12020_),
    .A2_N(_12022_),
    .B1(_11242_),
    .B2(_11917_),
    .Y(_12023_));
 sky130_fd_sc_hd__nor2_2 _28704_ (.A(_10813_),
    .B(_11917_),
    .Y(_12024_));
 sky130_fd_sc_hd__nand3_4 _28705_ (.A(_12022_),
    .B(_12020_),
    .C(_12024_),
    .Y(_12025_));
 sky130_fd_sc_hd__nand2_1 _28706_ (.A(_12023_),
    .B(_12025_),
    .Y(_12026_));
 sky130_fd_sc_hd__a21boi_1 _28707_ (.A1(_11928_),
    .A2(_11929_),
    .B1_N(_11927_),
    .Y(_12027_));
 sky130_fd_sc_hd__nand2_1 _28708_ (.A(_12026_),
    .B(_12027_),
    .Y(_12028_));
 sky130_fd_sc_hd__nand2_1 _28709_ (.A(_11931_),
    .B(_11927_),
    .Y(_12029_));
 sky130_fd_sc_hd__nand3_2 _28710_ (.A(_12029_),
    .B(_12023_),
    .C(_12025_),
    .Y(_12030_));
 sky130_fd_sc_hd__nand2_1 _28711_ (.A(_12028_),
    .B(_12030_),
    .Y(_12031_));
 sky130_fd_sc_hd__a21oi_1 _28712_ (.A1(_11941_),
    .A2(_11936_),
    .B1(_11935_),
    .Y(_12032_));
 sky130_fd_sc_hd__xor2_1 _28713_ (.A(_12031_),
    .B(_12032_),
    .X(_02674_));
 sky130_fd_sc_hd__clkbuf_4 _28714_ (.A(_11942_),
    .X(_12033_));
 sky130_fd_sc_hd__and2_1 _28715_ (.A(_11945_),
    .B(_11891_),
    .X(_12034_));
 sky130_fd_sc_hd__o21bai_4 _28716_ (.A1(_12033_),
    .A2(_11946_),
    .B1_N(_12034_),
    .Y(_12035_));
 sky130_fd_sc_hd__xor2_4 _28717_ (.A(_11361_),
    .B(_12035_),
    .X(_12036_));
 sky130_fd_sc_hd__xor2_1 _28718_ (.A(_11602_),
    .B(_12036_),
    .X(_12037_));
 sky130_vsdinv _28719_ (.A(_12037_),
    .Y(_12038_));
 sky130_fd_sc_hd__and2b_1 _28720_ (.A_N(_11949_),
    .B(_11993_),
    .X(_12039_));
 sky130_fd_sc_hd__o21bai_4 _28721_ (.A1(_11947_),
    .A2(_11994_),
    .B1_N(_12039_),
    .Y(_12040_));
 sky130_fd_sc_hd__buf_4 _28722_ (.A(_11943_),
    .X(_12041_));
 sky130_fd_sc_hd__buf_4 _28723_ (.A(_11892_),
    .X(_12042_));
 sky130_fd_sc_hd__nor2_1 _28724_ (.A(_11958_),
    .B(_11960_),
    .Y(_12043_));
 sky130_fd_sc_hd__o21bai_4 _28725_ (.A1(_11951_),
    .A2(_11961_),
    .B1_N(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__xor2_4 _28726_ (.A(_12042_),
    .B(_12044_),
    .X(_12045_));
 sky130_fd_sc_hd__xor2_4 _28727_ (.A(_12041_),
    .B(_12045_),
    .X(_12046_));
 sky130_fd_sc_hd__nor2_4 _28728_ (.A(_14006_),
    .B(_11953_),
    .Y(_12047_));
 sky130_fd_sc_hd__a21oi_4 _28729_ (.A1(_11957_),
    .A2(_11840_),
    .B1(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__a2bb2oi_4 _28730_ (.A1_N(_14006_),
    .A2_N(_11953_),
    .B1(_11744_),
    .B2(_11952_),
    .Y(_12049_));
 sky130_fd_sc_hd__xor2_4 _28731_ (.A(_12049_),
    .B(_11840_),
    .X(_12050_));
 sky130_fd_sc_hd__clkinv_16 _28732_ (.A(_12050_),
    .Y(_12051_));
 sky130_fd_sc_hd__nor2_1 _28733_ (.A(_11966_),
    .B(_11971_),
    .Y(_12052_));
 sky130_fd_sc_hd__o21bai_4 _28734_ (.A1(_11965_),
    .A2(_11972_),
    .B1_N(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__xor2_4 _28735_ (.A(_12051_),
    .B(_12053_),
    .X(_12054_));
 sky130_fd_sc_hd__xnor2_4 _28736_ (.A(_12048_),
    .B(_12054_),
    .Y(_12055_));
 sky130_fd_sc_hd__and2_1 _28737_ (.A(_11989_),
    .B(_11975_),
    .X(_12056_));
 sky130_fd_sc_hd__o21bai_4 _28738_ (.A1(_11973_),
    .A2(_11990_),
    .B1_N(_12056_),
    .Y(_12057_));
 sky130_fd_sc_hd__o21a_2 _28739_ (.A1(_11967_),
    .A2(_11970_),
    .B1(_11968_),
    .X(_12058_));
 sky130_fd_sc_hd__a2bb2oi_4 _28740_ (.A1_N(_14300_),
    .A2_N(_11977_),
    .B1(_11976_),
    .B2(_11978_),
    .Y(_12059_));
 sky130_fd_sc_hd__nand2_8 _28741_ (.A(_12780_),
    .B(net437),
    .Y(_12060_));
 sky130_fd_sc_hd__or4_4 _28742_ (.A(_13986_),
    .B(_13991_),
    .C(_14276_),
    .D(_14280_),
    .X(_12061_));
 sky130_fd_sc_hd__a22o_1 _28743_ (.A1(_11006_),
    .A2(_11138_),
    .B1(_07104_),
    .B2(_08596_),
    .X(_12062_));
 sky130_fd_sc_hd__nand2_2 _28744_ (.A(_12061_),
    .B(_12062_),
    .Y(_12063_));
 sky130_fd_sc_hd__xnor2_4 _28745_ (.A(_12060_),
    .B(_12063_),
    .Y(_12064_));
 sky130_fd_sc_hd__xnor2_4 _28746_ (.A(_12059_),
    .B(_12064_),
    .Y(_12065_));
 sky130_fd_sc_hd__xnor2_4 _28747_ (.A(_12058_),
    .B(_12065_),
    .Y(_12066_));
 sky130_fd_sc_hd__or2b_2 _28748_ (.A(_11987_),
    .B_N(_11982_),
    .X(_12067_));
 sky130_fd_sc_hd__o21ai_4 _28749_ (.A1(_11980_),
    .A2(_11988_),
    .B1(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__and2_2 _28750_ (.A(_07360_),
    .B(_08158_),
    .X(_12069_));
 sky130_fd_sc_hd__clkbuf_4 _28751_ (.A(_08397_),
    .X(_12070_));
 sky130_fd_sc_hd__nand3_4 _28752_ (.A(_12070_),
    .B(_11164_),
    .C(_07770_),
    .Y(_12071_));
 sky130_fd_sc_hd__a22o_2 _28753_ (.A1(_12070_),
    .A2(_07770_),
    .B1(_11164_),
    .B2(_08065_),
    .X(_12072_));
 sky130_fd_sc_hd__o21ai_4 _28754_ (.A1(_14293_),
    .A2(_12071_),
    .B1(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__xor2_4 _28755_ (.A(_12069_),
    .B(_12073_),
    .X(_12074_));
 sky130_fd_sc_hd__nand3b_2 _28756_ (.A_N(_11984_),
    .B(_08528_),
    .C(_14322_),
    .Y(_12075_));
 sky130_fd_sc_hd__o31ai_4 _28757_ (.A1(_13968_),
    .A2(_14311_),
    .A3(_11986_),
    .B1(_12075_),
    .Y(_12076_));
 sky130_fd_sc_hd__and2_2 _28758_ (.A(_07946_),
    .B(_10827_),
    .X(_12077_));
 sky130_fd_sc_hd__nand2_2 _28759_ (.A(_13962_),
    .B(_07467_),
    .Y(_12078_));
 sky130_fd_sc_hd__and2b_1 _28760_ (.A_N(_07198_),
    .B(_08526_),
    .X(_12079_));
 sky130_fd_sc_hd__xor2_4 _28761_ (.A(_12078_),
    .B(_12079_),
    .X(_12080_));
 sky130_fd_sc_hd__xor2_4 _28762_ (.A(_12077_),
    .B(_12080_),
    .X(_12081_));
 sky130_fd_sc_hd__xor2_4 _28763_ (.A(_12076_),
    .B(_12081_),
    .X(_12082_));
 sky130_fd_sc_hd__xor2_4 _28764_ (.A(_12074_),
    .B(_12082_),
    .X(_12083_));
 sky130_fd_sc_hd__xnor2_4 _28765_ (.A(_12068_),
    .B(_12083_),
    .Y(_12084_));
 sky130_fd_sc_hd__xor2_4 _28766_ (.A(_12066_),
    .B(_12084_),
    .X(_12085_));
 sky130_fd_sc_hd__xnor2_4 _28767_ (.A(_12057_),
    .B(_12085_),
    .Y(_12086_));
 sky130_fd_sc_hd__xor2_4 _28768_ (.A(_12055_),
    .B(_12086_),
    .X(_12087_));
 sky130_fd_sc_hd__and2b_1 _28769_ (.A_N(_11992_),
    .B(_11962_),
    .X(_12088_));
 sky130_fd_sc_hd__a21o_2 _28770_ (.A1(_11991_),
    .A2(_11964_),
    .B1(_12088_),
    .X(_12089_));
 sky130_fd_sc_hd__xnor2_4 _28771_ (.A(_12087_),
    .B(_12089_),
    .Y(_12090_));
 sky130_fd_sc_hd__xor2_4 _28772_ (.A(_12046_),
    .B(_12090_),
    .X(_12091_));
 sky130_fd_sc_hd__nor2_8 _28773_ (.A(_12040_),
    .B(_12091_),
    .Y(_12092_));
 sky130_fd_sc_hd__nand2_2 _28774_ (.A(_12091_),
    .B(_12040_),
    .Y(_12093_));
 sky130_fd_sc_hd__nor3b_4 _28775_ (.A(_12038_),
    .B(_12092_),
    .C_N(_12093_),
    .Y(_12094_));
 sky130_vsdinv _28776_ (.A(_12094_),
    .Y(_12095_));
 sky130_vsdinv _28777_ (.A(_12093_),
    .Y(_12096_));
 sky130_fd_sc_hd__o21bai_4 _28778_ (.A1(_12092_),
    .A2(_12096_),
    .B1_N(_12037_),
    .Y(_12097_));
 sky130_fd_sc_hd__o31ai_4 _28779_ (.A1(_12007_),
    .A2(_12008_),
    .A3(_11999_),
    .B1(_12000_),
    .Y(_12098_));
 sky130_fd_sc_hd__a21oi_4 _28780_ (.A1(_12095_),
    .A2(_12097_),
    .B1(_12098_),
    .Y(_12099_));
 sky130_fd_sc_hd__and3b_1 _28781_ (.A_N(_12094_),
    .B(_12097_),
    .C(_12098_),
    .X(_12100_));
 sky130_fd_sc_hd__buf_2 _28782_ (.A(_11473_),
    .X(_12101_));
 sky130_fd_sc_hd__o21ba_2 _28783_ (.A1(_12101_),
    .A2(_12004_),
    .B1_N(_12006_),
    .X(_12102_));
 sky130_fd_sc_hd__xor2_4 _28784_ (.A(_10812_),
    .B(_12102_),
    .X(_12103_));
 sky130_fd_sc_hd__o21bai_4 _28785_ (.A1(_12099_),
    .A2(_12100_),
    .B1_N(_12103_),
    .Y(_12104_));
 sky130_fd_sc_hd__nand3b_4 _28786_ (.A_N(_12094_),
    .B(_12097_),
    .C(_12098_),
    .Y(_12105_));
 sky130_fd_sc_hd__nand3b_4 _28787_ (.A_N(_12099_),
    .B(_12105_),
    .C(_12103_),
    .Y(_12106_));
 sky130_fd_sc_hd__nand2_2 _28788_ (.A(_12018_),
    .B(_12014_),
    .Y(_12107_));
 sky130_fd_sc_hd__a21oi_4 _28789_ (.A1(_12104_),
    .A2(_12106_),
    .B1(_12107_),
    .Y(_12108_));
 sky130_vsdinv _28790_ (.A(_12108_),
    .Y(_12109_));
 sky130_fd_sc_hd__nand3_4 _28791_ (.A(_12104_),
    .B(_12106_),
    .C(_12107_),
    .Y(_12110_));
 sky130_fd_sc_hd__nor2_1 _28792_ (.A(_11242_),
    .B(_12015_),
    .Y(_12111_));
 sky130_fd_sc_hd__a21oi_2 _28793_ (.A1(_12109_),
    .A2(_12110_),
    .B1(_12111_),
    .Y(_12112_));
 sky130_vsdinv _28794_ (.A(_12111_),
    .Y(_12113_));
 sky130_fd_sc_hd__nor3b_4 _28795_ (.A(_12113_),
    .B(_12108_),
    .C_N(_12110_),
    .Y(_12114_));
 sky130_vsdinv _28796_ (.A(_12114_),
    .Y(_12115_));
 sky130_fd_sc_hd__nand2_2 _28797_ (.A(_12025_),
    .B(_12020_),
    .Y(_12116_));
 sky130_fd_sc_hd__nand3b_4 _28798_ (.A_N(_12112_),
    .B(_12115_),
    .C(_12116_),
    .Y(_12117_));
 sky130_fd_sc_hd__o21bai_2 _28799_ (.A1(_12114_),
    .A2(_12112_),
    .B1_N(_12116_),
    .Y(_12118_));
 sky130_fd_sc_hd__nand2_4 _28800_ (.A(_12117_),
    .B(_12118_),
    .Y(_12119_));
 sky130_fd_sc_hd__nor3_2 _28801_ (.A(_11933_),
    .B(_11935_),
    .C(_12031_),
    .Y(_12120_));
 sky130_fd_sc_hd__nand2_1 _28802_ (.A(_11937_),
    .B(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__nand3_2 _28803_ (.A(_11508_),
    .B(_11507_),
    .C(_11626_),
    .Y(_12122_));
 sky130_fd_sc_hd__nor2_2 _28804_ (.A(_12121_),
    .B(_12122_),
    .Y(_12123_));
 sky130_fd_sc_hd__and2_1 _28805_ (.A(_12028_),
    .B(_12030_),
    .X(_12124_));
 sky130_fd_sc_hd__nand3_1 _28806_ (.A(_11936_),
    .B(_12124_),
    .C(_11940_),
    .Y(_12125_));
 sky130_fd_sc_hd__a21boi_1 _28807_ (.A1(_11935_),
    .A2(_12028_),
    .B1_N(_12030_),
    .Y(_12126_));
 sky130_fd_sc_hd__nand2_1 _28808_ (.A(_12125_),
    .B(_12126_),
    .Y(_12127_));
 sky130_fd_sc_hd__o21bai_2 _28809_ (.A1(_12121_),
    .A2(_11736_),
    .B1_N(_12127_),
    .Y(_12128_));
 sky130_fd_sc_hd__a21oi_4 _28810_ (.A1(_11269_),
    .A2(_12123_),
    .B1(_12128_),
    .Y(_12129_));
 sky130_fd_sc_hd__xor2_1 _28811_ (.A(_12119_),
    .B(_12129_),
    .X(_02675_));
 sky130_fd_sc_hd__buf_6 _28812_ (.A(_11361_),
    .X(_12130_));
 sky130_fd_sc_hd__and2_1 _28813_ (.A(_12035_),
    .B(_12130_),
    .X(_12131_));
 sky130_fd_sc_hd__a21oi_4 _28814_ (.A1(_12036_),
    .A2(net410),
    .B1(_12131_),
    .Y(_12132_));
 sky130_fd_sc_hd__xor2_4 _28815_ (.A(_10338_),
    .B(_12132_),
    .X(_12133_));
 sky130_vsdinv _28816_ (.A(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__nor2_2 _28817_ (.A(_12046_),
    .B(_12090_),
    .Y(_12135_));
 sky130_fd_sc_hd__and2_1 _28818_ (.A(_12053_),
    .B(_12050_),
    .X(_12136_));
 sky130_fd_sc_hd__o21bai_4 _28819_ (.A1(_12048_),
    .A2(_12054_),
    .B1_N(_12136_),
    .Y(_12137_));
 sky130_fd_sc_hd__xor2_4 _28820_ (.A(_12042_),
    .B(_12137_),
    .X(_12138_));
 sky130_fd_sc_hd__xor2_4 _28821_ (.A(_12041_),
    .B(_12138_),
    .X(_12139_));
 sky130_fd_sc_hd__and2_1 _28822_ (.A(_12085_),
    .B(_12057_),
    .X(_12140_));
 sky130_fd_sc_hd__o21bai_4 _28823_ (.A1(_12055_),
    .A2(_12086_),
    .B1_N(_12140_),
    .Y(_12141_));
 sky130_fd_sc_hd__nand2_1 _28824_ (.A(_11952_),
    .B(_11744_),
    .Y(_12142_));
 sky130_fd_sc_hd__a21oi_1 _28825_ (.A1(_11840_),
    .A2(_12142_),
    .B1(_12047_),
    .Y(_12143_));
 sky130_vsdinv _28826_ (.A(_12143_),
    .Y(_12144_));
 sky130_fd_sc_hd__nor2_1 _28827_ (.A(_12059_),
    .B(_12064_),
    .Y(_12145_));
 sky130_fd_sc_hd__o21bai_4 _28828_ (.A1(_12058_),
    .A2(_12065_),
    .B1_N(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__xor2_4 _28829_ (.A(_12051_),
    .B(_12146_),
    .X(_12147_));
 sky130_fd_sc_hd__xor2_4 _28830_ (.A(_12144_),
    .B(_12147_),
    .X(_12148_));
 sky130_fd_sc_hd__and2_1 _28831_ (.A(_12083_),
    .B(_12068_),
    .X(_12149_));
 sky130_fd_sc_hd__o21bai_4 _28832_ (.A1(_12066_),
    .A2(_12084_),
    .B1_N(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__o21a_2 _28833_ (.A1(_12060_),
    .A2(_12063_),
    .B1(_12061_),
    .X(_12151_));
 sky130_fd_sc_hd__a2bb2oi_4 _28834_ (.A1_N(_14294_),
    .A2_N(_12071_),
    .B1(_12069_),
    .B2(_12072_),
    .Y(_12152_));
 sky130_fd_sc_hd__nand2_2 _28835_ (.A(_11006_),
    .B(_08588_),
    .Y(_12153_));
 sky130_fd_sc_hd__nand2_8 _28836_ (.A(_12779_),
    .B(_07104_),
    .Y(_12154_));
 sky130_fd_sc_hd__xnor2_4 _28837_ (.A(_12153_),
    .B(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__xnor2_4 _28838_ (.A(_12060_),
    .B(_12155_),
    .Y(_12156_));
 sky130_fd_sc_hd__xnor2_4 _28839_ (.A(_12152_),
    .B(_12156_),
    .Y(_12157_));
 sky130_fd_sc_hd__xnor2_4 _28840_ (.A(_12151_),
    .B(_12157_),
    .Y(_12158_));
 sky130_fd_sc_hd__or2b_2 _28841_ (.A(_12081_),
    .B_N(_12076_),
    .X(_12159_));
 sky130_fd_sc_hd__o21ai_4 _28842_ (.A1(_12074_),
    .A2(_12082_),
    .B1(_12159_),
    .Y(_12160_));
 sky130_fd_sc_hd__and2_2 _28843_ (.A(_07360_),
    .B(_08482_),
    .X(_12161_));
 sky130_fd_sc_hd__nand3_4 _28844_ (.A(_13974_),
    .B(_13980_),
    .C(_08065_),
    .Y(_12162_));
 sky130_fd_sc_hd__a22o_2 _28845_ (.A1(_12070_),
    .A2(_08065_),
    .B1(_11164_),
    .B2(_08158_),
    .X(_12163_));
 sky130_fd_sc_hd__o21ai_4 _28846_ (.A1(_14286_),
    .A2(_12162_),
    .B1(_12163_),
    .Y(_12164_));
 sky130_fd_sc_hd__xor2_4 _28847_ (.A(_12161_),
    .B(_12164_),
    .X(_12165_));
 sky130_fd_sc_hd__nand3b_2 _28848_ (.A_N(_12078_),
    .B(_08528_),
    .C(_14316_),
    .Y(_12166_));
 sky130_fd_sc_hd__o31ai_4 _28849_ (.A1(_13968_),
    .A2(_14305_),
    .A3(_12080_),
    .B1(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__and2_2 _28850_ (.A(_07946_),
    .B(_10829_),
    .X(_12168_));
 sky130_fd_sc_hd__nand2_2 _28851_ (.A(_13962_),
    .B(_07775_),
    .Y(_12169_));
 sky130_fd_sc_hd__and2b_1 _28852_ (.A_N(_07467_),
    .B(_09169_),
    .X(_12170_));
 sky130_fd_sc_hd__xor2_4 _28853_ (.A(_12169_),
    .B(_12170_),
    .X(_12171_));
 sky130_fd_sc_hd__xor2_4 _28854_ (.A(_12168_),
    .B(_12171_),
    .X(_12172_));
 sky130_fd_sc_hd__xor2_4 _28855_ (.A(_12167_),
    .B(_12172_),
    .X(_12173_));
 sky130_fd_sc_hd__xor2_4 _28856_ (.A(_12165_),
    .B(_12173_),
    .X(_12174_));
 sky130_fd_sc_hd__xnor2_4 _28857_ (.A(_12160_),
    .B(_12174_),
    .Y(_12175_));
 sky130_fd_sc_hd__xor2_4 _28858_ (.A(_12158_),
    .B(_12175_),
    .X(_12176_));
 sky130_fd_sc_hd__xnor2_4 _28859_ (.A(_12150_),
    .B(_12176_),
    .Y(_12177_));
 sky130_fd_sc_hd__xor2_4 _28860_ (.A(_12148_),
    .B(_12177_),
    .X(_12178_));
 sky130_fd_sc_hd__xnor2_4 _28861_ (.A(_12141_),
    .B(_12178_),
    .Y(_12179_));
 sky130_fd_sc_hd__xor2_4 _28862_ (.A(_12139_),
    .B(_12179_),
    .X(_12180_));
 sky130_fd_sc_hd__a211oi_4 _28863_ (.A1(_12087_),
    .A2(_12089_),
    .B1(_12135_),
    .C1(_12180_),
    .Y(_12181_));
 sky130_fd_sc_hd__a21o_1 _28864_ (.A1(_12087_),
    .A2(_12089_),
    .B1(_12135_),
    .X(_12182_));
 sky130_fd_sc_hd__nand2_4 _28865_ (.A(_12182_),
    .B(_12180_),
    .Y(_12183_));
 sky130_vsdinv _28866_ (.A(_12183_),
    .Y(_12184_));
 sky130_fd_sc_hd__nand2_1 _28867_ (.A(_12044_),
    .B(_12002_),
    .Y(_12185_));
 sky130_fd_sc_hd__o21a_2 _28868_ (.A1(_12033_),
    .A2(_12045_),
    .B1(_12185_),
    .X(_12186_));
 sky130_fd_sc_hd__xor2_4 _28869_ (.A(_11489_),
    .B(_12186_),
    .X(_12187_));
 sky130_fd_sc_hd__xor2_4 _28870_ (.A(_11602_),
    .B(_12187_),
    .X(_12188_));
 sky130_fd_sc_hd__o21bai_4 _28871_ (.A1(_12181_),
    .A2(_12184_),
    .B1_N(_12188_),
    .Y(_12189_));
 sky130_fd_sc_hd__nand3b_4 _28872_ (.A_N(_12181_),
    .B(_12183_),
    .C(_12188_),
    .Y(_12190_));
 sky130_fd_sc_hd__o21ai_4 _28873_ (.A1(_12038_),
    .A2(_12092_),
    .B1(_12093_),
    .Y(_12191_));
 sky130_fd_sc_hd__a21oi_4 _28874_ (.A1(_12189_),
    .A2(_12190_),
    .B1(_12191_),
    .Y(_12192_));
 sky130_fd_sc_hd__nand3_4 _28875_ (.A(_12189_),
    .B(_12191_),
    .C(_12190_),
    .Y(_12193_));
 sky130_fd_sc_hd__nor3b_4 _28876_ (.A(_12134_),
    .B(_12192_),
    .C_N(_12193_),
    .Y(_12194_));
 sky130_vsdinv _28877_ (.A(_12192_),
    .Y(_12195_));
 sky130_fd_sc_hd__a21oi_4 _28878_ (.A1(_12195_),
    .A2(_12193_),
    .B1(_12133_),
    .Y(_12196_));
 sky130_fd_sc_hd__a211o_2 _28879_ (.A1(_12106_),
    .A2(_12105_),
    .B1(_12194_),
    .C1(_12196_),
    .X(_12197_));
 sky130_fd_sc_hd__o211ai_4 _28880_ (.A1(_12194_),
    .A2(_12196_),
    .B1(_12105_),
    .C1(_12106_),
    .Y(_12198_));
 sky130_fd_sc_hd__nor2_2 _28881_ (.A(_11243_),
    .B(_12102_),
    .Y(_12199_));
 sky130_fd_sc_hd__a21o_1 _28882_ (.A1(_12197_),
    .A2(_12198_),
    .B1(_12199_),
    .X(_12200_));
 sky130_fd_sc_hd__nand3_4 _28883_ (.A(_12197_),
    .B(_12198_),
    .C(_12199_),
    .Y(_12201_));
 sky130_fd_sc_hd__o21ai_4 _28884_ (.A1(_12113_),
    .A2(_12108_),
    .B1(_12110_),
    .Y(_12202_));
 sky130_fd_sc_hd__a21oi_4 _28885_ (.A1(_12200_),
    .A2(_12201_),
    .B1(_12202_),
    .Y(_12203_));
 sky130_fd_sc_hd__nand3_4 _28886_ (.A(_12200_),
    .B(_12201_),
    .C(_12202_),
    .Y(_12204_));
 sky130_fd_sc_hd__or2b_2 _28887_ (.A(_12203_),
    .B_N(_12204_),
    .X(_12205_));
 sky130_fd_sc_hd__o21a_1 _28888_ (.A1(_12119_),
    .A2(_12129_),
    .B1(_12117_),
    .X(_12206_));
 sky130_fd_sc_hd__xor2_1 _28889_ (.A(_12205_),
    .B(_12206_),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_1 _28890_ (.A(_12137_),
    .B(_11891_),
    .Y(_12207_));
 sky130_fd_sc_hd__o21a_2 _28891_ (.A1(_11942_),
    .A2(_12138_),
    .B1(_12207_),
    .X(_12208_));
 sky130_fd_sc_hd__xor2_4 _28892_ (.A(_11361_),
    .B(_12208_),
    .X(_12209_));
 sky130_fd_sc_hd__xor2_4 _28893_ (.A(_11473_),
    .B(_12209_),
    .X(_12210_));
 sky130_vsdinv _28894_ (.A(_12210_),
    .Y(_12211_));
 sky130_fd_sc_hd__buf_4 _28895_ (.A(_12143_),
    .X(_12212_));
 sky130_fd_sc_hd__clkbuf_4 _28896_ (.A(_12050_),
    .X(_12213_));
 sky130_fd_sc_hd__and2_1 _28897_ (.A(_12146_),
    .B(_12213_),
    .X(_12214_));
 sky130_fd_sc_hd__o21bai_4 _28898_ (.A1(_12212_),
    .A2(_12147_),
    .B1_N(_12214_),
    .Y(_12215_));
 sky130_fd_sc_hd__xor2_4 _28899_ (.A(net411),
    .B(_12215_),
    .X(_12216_));
 sky130_fd_sc_hd__xor2_4 _28900_ (.A(net412),
    .B(_12216_),
    .X(_12217_));
 sky130_fd_sc_hd__and2_1 _28901_ (.A(_12176_),
    .B(_12150_),
    .X(_12218_));
 sky130_fd_sc_hd__o21bai_4 _28902_ (.A1(_12148_),
    .A2(_12177_),
    .B1_N(_12218_),
    .Y(_12219_));
 sky130_fd_sc_hd__nor2_1 _28903_ (.A(_12152_),
    .B(_12156_),
    .Y(_12220_));
 sky130_fd_sc_hd__o21bai_4 _28904_ (.A1(_12151_),
    .A2(_12157_),
    .B1_N(_12220_),
    .Y(_12221_));
 sky130_fd_sc_hd__xor2_4 _28905_ (.A(_12051_),
    .B(_12221_),
    .X(_12222_));
 sky130_fd_sc_hd__xor2_4 _28906_ (.A(_12144_),
    .B(_12222_),
    .X(_12223_));
 sky130_fd_sc_hd__and2_1 _28907_ (.A(_12174_),
    .B(_12160_),
    .X(_12224_));
 sky130_fd_sc_hd__o21bai_4 _28908_ (.A1(_12158_),
    .A2(_12175_),
    .B1_N(_12224_),
    .Y(_12225_));
 sky130_fd_sc_hd__nand3b_1 _28909_ (.A_N(_12154_),
    .B(_11006_),
    .C(_08589_),
    .Y(_12226_));
 sky130_fd_sc_hd__o21a_2 _28910_ (.A1(_12060_),
    .A2(_12155_),
    .B1(_12226_),
    .X(_12227_));
 sky130_fd_sc_hd__o2bb2ai_4 _28911_ (.A1_N(_12163_),
    .A2_N(_12161_),
    .B1(_14287_),
    .B2(_12162_),
    .Y(_12228_));
 sky130_fd_sc_hd__nand2_2 _28912_ (.A(_09468_),
    .B(_11006_),
    .Y(_12229_));
 sky130_fd_sc_hd__xnor2_4 _28913_ (.A(_12154_),
    .B(_12229_),
    .Y(_12230_));
 sky130_fd_sc_hd__xor2_4 _28914_ (.A(_12060_),
    .B(_12230_),
    .X(_12231_));
 sky130_fd_sc_hd__xnor2_4 _28915_ (.A(_12228_),
    .B(_12231_),
    .Y(_12232_));
 sky130_fd_sc_hd__xnor2_4 _28916_ (.A(_12227_),
    .B(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__or2b_2 _28917_ (.A(_12172_),
    .B_N(_12167_),
    .X(_12234_));
 sky130_fd_sc_hd__o21ai_4 _28918_ (.A1(_12165_),
    .A2(_12173_),
    .B1(_12234_),
    .Y(_12235_));
 sky130_fd_sc_hd__and2_2 _28919_ (.A(_07360_),
    .B(_08589_),
    .X(_12236_));
 sky130_fd_sc_hd__nand3_4 _28920_ (.A(_13974_),
    .B(_13980_),
    .C(_08158_),
    .Y(_12237_));
 sky130_fd_sc_hd__a22o_2 _28921_ (.A1(_12070_),
    .A2(_08158_),
    .B1(_13980_),
    .B2(_08481_),
    .X(_12238_));
 sky130_fd_sc_hd__o21ai_4 _28922_ (.A1(_14281_),
    .A2(_12237_),
    .B1(_12238_),
    .Y(_12239_));
 sky130_fd_sc_hd__xor2_4 _28923_ (.A(_12236_),
    .B(_12239_),
    .X(_12240_));
 sky130_fd_sc_hd__nand3b_2 _28924_ (.A_N(_12169_),
    .B(_08528_),
    .C(_14310_),
    .Y(_12241_));
 sky130_fd_sc_hd__o31ai_4 _28925_ (.A1(_13969_),
    .A2(_14299_),
    .A3(_12171_),
    .B1(_12241_),
    .Y(_12242_));
 sky130_fd_sc_hd__and2_2 _28926_ (.A(_08244_),
    .B(_10825_),
    .X(_12243_));
 sky130_fd_sc_hd__nand2_2 _28927_ (.A(_13962_),
    .B(_07769_),
    .Y(_12244_));
 sky130_fd_sc_hd__and2b_2 _28928_ (.A_N(_07569_),
    .B(_09169_),
    .X(_12245_));
 sky130_fd_sc_hd__xor2_4 _28929_ (.A(_12244_),
    .B(_12245_),
    .X(_12246_));
 sky130_fd_sc_hd__xor2_4 _28930_ (.A(_12243_),
    .B(_12246_),
    .X(_12247_));
 sky130_fd_sc_hd__xor2_4 _28931_ (.A(_12242_),
    .B(_12247_),
    .X(_12248_));
 sky130_fd_sc_hd__xor2_4 _28932_ (.A(_12240_),
    .B(_12248_),
    .X(_12249_));
 sky130_fd_sc_hd__xnor2_4 _28933_ (.A(_12235_),
    .B(_12249_),
    .Y(_12250_));
 sky130_fd_sc_hd__xor2_4 _28934_ (.A(_12233_),
    .B(_12250_),
    .X(_12251_));
 sky130_fd_sc_hd__xnor2_4 _28935_ (.A(_12225_),
    .B(_12251_),
    .Y(_12252_));
 sky130_fd_sc_hd__xor2_4 _28936_ (.A(_12223_),
    .B(_12252_),
    .X(_12253_));
 sky130_fd_sc_hd__xnor2_4 _28937_ (.A(_12219_),
    .B(_12253_),
    .Y(_12254_));
 sky130_fd_sc_hd__xor2_4 _28938_ (.A(_12217_),
    .B(_12254_),
    .X(_12255_));
 sky130_fd_sc_hd__nor2_1 _28939_ (.A(_12139_),
    .B(_12179_),
    .Y(_12256_));
 sky130_fd_sc_hd__a21o_2 _28940_ (.A1(_12178_),
    .A2(_12141_),
    .B1(_12256_),
    .X(_12257_));
 sky130_fd_sc_hd__nor2_4 _28941_ (.A(_12255_),
    .B(_12257_),
    .Y(_12258_));
 sky130_fd_sc_hd__nand2_4 _28942_ (.A(_12257_),
    .B(_12255_),
    .Y(_12259_));
 sky130_fd_sc_hd__nor3b_4 _28943_ (.A(_12211_),
    .B(_12258_),
    .C_N(_12259_),
    .Y(_12260_));
 sky130_vsdinv _28944_ (.A(_12258_),
    .Y(_12261_));
 sky130_fd_sc_hd__a21oi_4 _28945_ (.A1(_12261_),
    .A2(_12259_),
    .B1(_12210_),
    .Y(_12262_));
 sky130_fd_sc_hd__a211oi_4 _28946_ (.A1(_12190_),
    .A2(_12183_),
    .B1(_12260_),
    .C1(_12262_),
    .Y(_12263_));
 sky130_fd_sc_hd__o211a_2 _28947_ (.A1(_12260_),
    .A2(_12262_),
    .B1(_12183_),
    .C1(_12190_),
    .X(_12264_));
 sky130_fd_sc_hd__nor2_2 _28948_ (.A(_11489_),
    .B(_12186_),
    .Y(_12265_));
 sky130_fd_sc_hd__a21oi_4 _28949_ (.A1(_12187_),
    .A2(net410),
    .B1(_12265_),
    .Y(_12266_));
 sky130_fd_sc_hd__xor2_1 _28950_ (.A(_10338_),
    .B(_12266_),
    .X(_12267_));
 sky130_vsdinv _28951_ (.A(_12267_),
    .Y(_12268_));
 sky130_fd_sc_hd__o21a_1 _28952_ (.A1(_12263_),
    .A2(_12264_),
    .B1(_12268_),
    .X(_12269_));
 sky130_fd_sc_hd__a211o_1 _28953_ (.A1(_12190_),
    .A2(_12183_),
    .B1(_12260_),
    .C1(_12262_),
    .X(_12270_));
 sky130_fd_sc_hd__nor3b_4 _28954_ (.A(_12268_),
    .B(_12264_),
    .C_N(_12270_),
    .Y(_12271_));
 sky130_vsdinv _28955_ (.A(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__o21ai_2 _28956_ (.A1(_12134_),
    .A2(_12192_),
    .B1(_12193_),
    .Y(_12273_));
 sky130_fd_sc_hd__nand3b_4 _28957_ (.A_N(_12269_),
    .B(_12272_),
    .C(_12273_),
    .Y(_12274_));
 sky130_fd_sc_hd__o21bai_4 _28958_ (.A1(_12269_),
    .A2(_12271_),
    .B1_N(_12273_),
    .Y(_12275_));
 sky130_fd_sc_hd__nor2_8 _28959_ (.A(_11243_),
    .B(_12132_),
    .Y(_12276_));
 sky130_fd_sc_hd__a21oi_1 _28960_ (.A1(_12274_),
    .A2(_12275_),
    .B1(_12276_),
    .Y(_12277_));
 sky130_vsdinv _28961_ (.A(_12277_),
    .Y(_12278_));
 sky130_fd_sc_hd__nand3_4 _28962_ (.A(_12274_),
    .B(_12276_),
    .C(_12275_),
    .Y(_12279_));
 sky130_fd_sc_hd__nand2_2 _28963_ (.A(_12201_),
    .B(_12197_),
    .Y(_12280_));
 sky130_fd_sc_hd__a21o_1 _28964_ (.A1(_12278_),
    .A2(_12279_),
    .B1(_12280_),
    .X(_12281_));
 sky130_fd_sc_hd__nand3_4 _28965_ (.A(_12278_),
    .B(_12280_),
    .C(_12279_),
    .Y(_12282_));
 sky130_fd_sc_hd__nand2_1 _28966_ (.A(_12281_),
    .B(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__a21oi_4 _28967_ (.A1(_12117_),
    .A2(_12204_),
    .B1(_12203_),
    .Y(_12284_));
 sky130_fd_sc_hd__nor3_4 _28968_ (.A(_12119_),
    .B(_12205_),
    .C(_12129_),
    .Y(_12285_));
 sky130_fd_sc_hd__nor2_2 _28969_ (.A(_12284_),
    .B(_12285_),
    .Y(_12286_));
 sky130_fd_sc_hd__xor2_1 _28970_ (.A(_12283_),
    .B(_12286_),
    .X(_02677_));
 sky130_vsdinv _28971_ (.A(_12282_),
    .Y(_12287_));
 sky130_fd_sc_hd__a21oi_1 _28972_ (.A1(_12278_),
    .A2(_12279_),
    .B1(_12280_),
    .Y(_12288_));
 sky130_fd_sc_hd__nor2_2 _28973_ (.A(_12288_),
    .B(_12287_),
    .Y(_12289_));
 sky130_fd_sc_hd__o21a_1 _28974_ (.A1(_12284_),
    .A2(_12285_),
    .B1(_12289_),
    .X(_12290_));
 sky130_fd_sc_hd__nand2_1 _28975_ (.A(_12215_),
    .B(_12002_),
    .Y(_12291_));
 sky130_fd_sc_hd__o21a_1 _28976_ (.A1(_12033_),
    .A2(_12216_),
    .B1(_12291_),
    .X(_12292_));
 sky130_fd_sc_hd__xor2_2 _28977_ (.A(_11361_),
    .B(_12292_),
    .X(_12293_));
 sky130_fd_sc_hd__xor2_1 _28978_ (.A(_11473_),
    .B(_12293_),
    .X(_12294_));
 sky130_vsdinv _28979_ (.A(_12294_),
    .Y(_12295_));
 sky130_fd_sc_hd__and2_1 _28980_ (.A(_12253_),
    .B(_12219_),
    .X(_12296_));
 sky130_fd_sc_hd__o21bai_2 _28981_ (.A1(_12217_),
    .A2(_12254_),
    .B1_N(_12296_),
    .Y(_12297_));
 sky130_fd_sc_hd__and2_1 _28982_ (.A(_12221_),
    .B(_12213_),
    .X(_12298_));
 sky130_fd_sc_hd__o21bai_4 _28983_ (.A1(_12212_),
    .A2(_12222_),
    .B1_N(_12298_),
    .Y(_12299_));
 sky130_fd_sc_hd__xor2_4 _28984_ (.A(net411),
    .B(_12299_),
    .X(_12300_));
 sky130_fd_sc_hd__xor2_4 _28985_ (.A(net412),
    .B(_12300_),
    .X(_12301_));
 sky130_fd_sc_hd__and2_1 _28986_ (.A(_12251_),
    .B(_12225_),
    .X(_12302_));
 sky130_fd_sc_hd__o21bai_2 _28987_ (.A1(_12223_),
    .A2(_12252_),
    .B1_N(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__and2_1 _28988_ (.A(_12231_),
    .B(_12228_),
    .X(_12304_));
 sky130_fd_sc_hd__o21bai_4 _28989_ (.A1(_12227_),
    .A2(_12232_),
    .B1_N(_12304_),
    .Y(_12305_));
 sky130_fd_sc_hd__xor2_4 _28990_ (.A(_12051_),
    .B(_12305_),
    .X(_12306_));
 sky130_fd_sc_hd__xor2_4 _28991_ (.A(_12144_),
    .B(_12306_),
    .X(_12307_));
 sky130_fd_sc_hd__and2_1 _28992_ (.A(_12249_),
    .B(_12235_),
    .X(_12308_));
 sky130_fd_sc_hd__o21bai_4 _28993_ (.A1(_12233_),
    .A2(_12250_),
    .B1_N(_12308_),
    .Y(_12309_));
 sky130_fd_sc_hd__o22a_4 _28994_ (.A1(_13986_),
    .A2(_12154_),
    .B1(_12060_),
    .B2(_12230_),
    .X(_12310_));
 sky130_fd_sc_hd__o2bb2ai_4 _28995_ (.A1_N(_12238_),
    .A2_N(_12236_),
    .B1(_14281_),
    .B2(_12237_),
    .Y(_12311_));
 sky130_fd_sc_hd__xnor2_4 _28996_ (.A(_12311_),
    .B(_12231_),
    .Y(_12312_));
 sky130_fd_sc_hd__xnor2_4 _28997_ (.A(_12310_),
    .B(_12312_),
    .Y(_12313_));
 sky130_fd_sc_hd__or2b_1 _28998_ (.A(_12247_),
    .B_N(_12242_),
    .X(_12314_));
 sky130_fd_sc_hd__o21ai_4 _28999_ (.A1(_12240_),
    .A2(_12248_),
    .B1(_12314_),
    .Y(_12315_));
 sky130_fd_sc_hd__and2_1 _29000_ (.A(_09468_),
    .B(_11162_),
    .X(_12316_));
 sky130_fd_sc_hd__buf_6 _29001_ (.A(_12316_),
    .X(_12317_));
 sky130_fd_sc_hd__nand3_4 _29002_ (.A(_13974_),
    .B(_13980_),
    .C(_08482_),
    .Y(_12318_));
 sky130_fd_sc_hd__a22o_2 _29003_ (.A1(_12070_),
    .A2(_08481_),
    .B1(_13980_),
    .B2(_08588_),
    .X(_12319_));
 sky130_fd_sc_hd__o21ai_4 _29004_ (.A1(_14276_),
    .A2(_12318_),
    .B1(_12319_),
    .Y(_12320_));
 sky130_fd_sc_hd__xor2_4 _29005_ (.A(_12317_),
    .B(_12320_),
    .X(_12321_));
 sky130_fd_sc_hd__nand3b_2 _29006_ (.A_N(_12244_),
    .B(_08528_),
    .C(_14305_),
    .Y(_12322_));
 sky130_fd_sc_hd__o31ai_4 _29007_ (.A1(_13969_),
    .A2(_14293_),
    .A3(_12246_),
    .B1(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__and2_2 _29008_ (.A(_08244_),
    .B(_08489_),
    .X(_12324_));
 sky130_fd_sc_hd__nand2_2 _29009_ (.A(_13963_),
    .B(_08064_),
    .Y(_12325_));
 sky130_fd_sc_hd__and2b_2 _29010_ (.A_N(_08070_),
    .B(_09876_),
    .X(_12326_));
 sky130_fd_sc_hd__xor2_4 _29011_ (.A(_12325_),
    .B(_12326_),
    .X(_12327_));
 sky130_fd_sc_hd__xor2_4 _29012_ (.A(_12324_),
    .B(_12327_),
    .X(_12328_));
 sky130_fd_sc_hd__xor2_4 _29013_ (.A(_12323_),
    .B(_12328_),
    .X(_12329_));
 sky130_fd_sc_hd__xor2_4 _29014_ (.A(_12321_),
    .B(_12329_),
    .X(_12330_));
 sky130_fd_sc_hd__xnor2_4 _29015_ (.A(_12315_),
    .B(_12330_),
    .Y(_12331_));
 sky130_fd_sc_hd__xor2_4 _29016_ (.A(_12313_),
    .B(_12331_),
    .X(_12332_));
 sky130_fd_sc_hd__xnor2_4 _29017_ (.A(_12309_),
    .B(_12332_),
    .Y(_12333_));
 sky130_fd_sc_hd__xor2_4 _29018_ (.A(_12307_),
    .B(_12333_),
    .X(_12334_));
 sky130_fd_sc_hd__xnor2_2 _29019_ (.A(_12303_),
    .B(_12334_),
    .Y(_12335_));
 sky130_fd_sc_hd__xor2_2 _29020_ (.A(_12301_),
    .B(_12335_),
    .X(_12336_));
 sky130_fd_sc_hd__xnor2_1 _29021_ (.A(_12297_),
    .B(_12336_),
    .Y(_12337_));
 sky130_fd_sc_hd__nor2_2 _29022_ (.A(_12295_),
    .B(_12337_),
    .Y(_12338_));
 sky130_vsdinv _29023_ (.A(_12338_),
    .Y(_12339_));
 sky130_fd_sc_hd__nand2_2 _29024_ (.A(_12337_),
    .B(_12295_),
    .Y(_12340_));
 sky130_fd_sc_hd__o21ai_4 _29025_ (.A1(_12211_),
    .A2(_12258_),
    .B1(_12259_),
    .Y(_12341_));
 sky130_fd_sc_hd__a21oi_4 _29026_ (.A1(_12339_),
    .A2(_12340_),
    .B1(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__and3b_1 _29027_ (.A_N(_12338_),
    .B(_12340_),
    .C(_12341_),
    .X(_12343_));
 sky130_fd_sc_hd__nor2_1 _29028_ (.A(_11489_),
    .B(_12208_),
    .Y(_12344_));
 sky130_fd_sc_hd__o21ba_2 _29029_ (.A1(_12101_),
    .A2(_12209_),
    .B1_N(_12344_),
    .X(_12345_));
 sky130_fd_sc_hd__xor2_1 _29030_ (.A(_10338_),
    .B(_12345_),
    .X(_12346_));
 sky130_vsdinv _29031_ (.A(_12346_),
    .Y(_12347_));
 sky130_fd_sc_hd__o21a_1 _29032_ (.A1(_12342_),
    .A2(_12343_),
    .B1(_12347_),
    .X(_12348_));
 sky130_fd_sc_hd__nand3b_4 _29033_ (.A_N(_12338_),
    .B(_12340_),
    .C(_12341_),
    .Y(_12349_));
 sky130_fd_sc_hd__nor3b_4 _29034_ (.A(_12347_),
    .B(_12342_),
    .C_N(_12349_),
    .Y(_12350_));
 sky130_vsdinv _29035_ (.A(_12350_),
    .Y(_12351_));
 sky130_fd_sc_hd__o21ai_2 _29036_ (.A1(_12268_),
    .A2(_12264_),
    .B1(_12270_),
    .Y(_12352_));
 sky130_fd_sc_hd__nand3b_4 _29037_ (.A_N(_12348_),
    .B(_12351_),
    .C(_12352_),
    .Y(_12353_));
 sky130_fd_sc_hd__o21bai_2 _29038_ (.A1(_12350_),
    .A2(_12348_),
    .B1_N(_12352_),
    .Y(_12354_));
 sky130_fd_sc_hd__nor2_2 _29039_ (.A(_11615_),
    .B(_12266_),
    .Y(_12355_));
 sky130_fd_sc_hd__a21oi_4 _29040_ (.A1(_12353_),
    .A2(_12354_),
    .B1(_12355_),
    .Y(_12356_));
 sky130_fd_sc_hd__nand3_1 _29041_ (.A(_12353_),
    .B(_12355_),
    .C(_12354_),
    .Y(_12357_));
 sky130_vsdinv _29042_ (.A(_12357_),
    .Y(_12358_));
 sky130_fd_sc_hd__a21boi_4 _29043_ (.A1(_12275_),
    .A2(_12276_),
    .B1_N(_12274_),
    .Y(_12359_));
 sky130_fd_sc_hd__o21a_1 _29044_ (.A1(_12356_),
    .A2(_12358_),
    .B1(_12359_),
    .X(_12360_));
 sky130_fd_sc_hd__nor3_4 _29045_ (.A(_12356_),
    .B(_12358_),
    .C(_12359_),
    .Y(_12361_));
 sky130_fd_sc_hd__nor2_4 _29046_ (.A(_12360_),
    .B(_12361_),
    .Y(_12362_));
 sky130_fd_sc_hd__o21bai_1 _29047_ (.A1(_12287_),
    .A2(_12290_),
    .B1_N(_12362_),
    .Y(_12363_));
 sky130_fd_sc_hd__o211ai_1 _29048_ (.A1(_12283_),
    .A2(_12286_),
    .B1(_12282_),
    .C1(_12362_),
    .Y(_12364_));
 sky130_fd_sc_hd__nand2_1 _29049_ (.A(_12363_),
    .B(_12364_),
    .Y(_02678_));
 sky130_fd_sc_hd__nor2_1 _29050_ (.A(_11489_),
    .B(_12292_),
    .Y(_12365_));
 sky130_fd_sc_hd__o21ba_2 _29051_ (.A1(_12101_),
    .A2(_12293_),
    .B1_N(_12365_),
    .X(_12366_));
 sky130_fd_sc_hd__xor2_1 _29052_ (.A(_10812_),
    .B(_12366_),
    .X(_12367_));
 sky130_vsdinv _29053_ (.A(_12367_),
    .Y(_12368_));
 sky130_fd_sc_hd__a21o_1 _29054_ (.A1(_12336_),
    .A2(_12297_),
    .B1(_12338_),
    .X(_12369_));
 sky130_fd_sc_hd__nand2_1 _29055_ (.A(_12299_),
    .B(_12002_),
    .Y(_12370_));
 sky130_fd_sc_hd__o21a_2 _29056_ (.A1(_12033_),
    .A2(_12300_),
    .B1(_12370_),
    .X(_12371_));
 sky130_fd_sc_hd__xor2_4 _29057_ (.A(_12130_),
    .B(_12371_),
    .X(_12372_));
 sky130_fd_sc_hd__xor2_4 _29058_ (.A(net410),
    .B(_12372_),
    .X(_12373_));
 sky130_fd_sc_hd__and2_1 _29059_ (.A(_12305_),
    .B(_12213_),
    .X(_12374_));
 sky130_fd_sc_hd__o21bai_4 _29060_ (.A1(_12212_),
    .A2(_12306_),
    .B1_N(_12374_),
    .Y(_12375_));
 sky130_fd_sc_hd__xor2_4 _29061_ (.A(net411),
    .B(_12375_),
    .X(_12376_));
 sky130_fd_sc_hd__xor2_4 _29062_ (.A(net412),
    .B(_12376_),
    .X(_12377_));
 sky130_fd_sc_hd__and2_1 _29063_ (.A(_12332_),
    .B(_12309_),
    .X(_12378_));
 sky130_fd_sc_hd__o21bai_4 _29064_ (.A1(_12307_),
    .A2(_12333_),
    .B1_N(_12378_),
    .Y(_12379_));
 sky130_fd_sc_hd__buf_6 _29065_ (.A(_12310_),
    .X(_12380_));
 sky130_fd_sc_hd__buf_4 _29066_ (.A(_12231_),
    .X(_12381_));
 sky130_fd_sc_hd__and2_1 _29067_ (.A(_12381_),
    .B(_12311_),
    .X(_12382_));
 sky130_fd_sc_hd__o21bai_4 _29068_ (.A1(_12380_),
    .A2(_12312_),
    .B1_N(_12382_),
    .Y(_12383_));
 sky130_fd_sc_hd__xor2_4 _29069_ (.A(_12051_),
    .B(_12383_),
    .X(_12384_));
 sky130_fd_sc_hd__xor2_4 _29070_ (.A(_12144_),
    .B(_12384_),
    .X(_12385_));
 sky130_fd_sc_hd__and2_1 _29071_ (.A(_12330_),
    .B(_12315_),
    .X(_12386_));
 sky130_fd_sc_hd__o21bai_4 _29072_ (.A1(_12313_),
    .A2(_12331_),
    .B1_N(_12386_),
    .Y(_12387_));
 sky130_fd_sc_hd__o2bb2ai_4 _29073_ (.A1_N(_12319_),
    .A2_N(_12317_),
    .B1(_14277_),
    .B2(_12318_),
    .Y(_12388_));
 sky130_fd_sc_hd__xnor2_4 _29074_ (.A(_12388_),
    .B(_12381_),
    .Y(_12389_));
 sky130_fd_sc_hd__xnor2_4 _29075_ (.A(_12380_),
    .B(_12389_),
    .Y(_12390_));
 sky130_fd_sc_hd__or2b_2 _29076_ (.A(_12328_),
    .B_N(_12323_),
    .X(_12391_));
 sky130_fd_sc_hd__o21ai_4 _29077_ (.A1(_12321_),
    .A2(_12329_),
    .B1(_12391_),
    .Y(_12392_));
 sky130_fd_sc_hd__nand2_2 _29078_ (.A(_13974_),
    .B(_08589_),
    .Y(_12393_));
 sky130_fd_sc_hd__nand2_8 _29079_ (.A(_09468_),
    .B(_11164_),
    .Y(_12394_));
 sky130_fd_sc_hd__xnor2_4 _29080_ (.A(_12393_),
    .B(_12394_),
    .Y(_12395_));
 sky130_fd_sc_hd__xor2_4 _29081_ (.A(_12317_),
    .B(_12395_),
    .X(_12396_));
 sky130_fd_sc_hd__nand3b_2 _29082_ (.A_N(_12325_),
    .B(_08529_),
    .C(_14300_),
    .Y(_12397_));
 sky130_fd_sc_hd__o31ai_4 _29083_ (.A1(_13969_),
    .A2(_14287_),
    .A3(_12327_),
    .B1(_12397_),
    .Y(_12398_));
 sky130_fd_sc_hd__and2_2 _29084_ (.A(_08244_),
    .B(_08481_),
    .X(_12399_));
 sky130_fd_sc_hd__nand2_2 _29085_ (.A(_13963_),
    .B(_08489_),
    .Y(_12400_));
 sky130_fd_sc_hd__and2b_1 _29086_ (.A_N(_10825_),
    .B(_08527_),
    .X(_12401_));
 sky130_fd_sc_hd__xor2_4 _29087_ (.A(_12400_),
    .B(_12401_),
    .X(_12402_));
 sky130_fd_sc_hd__xor2_4 _29088_ (.A(_12399_),
    .B(_12402_),
    .X(_12403_));
 sky130_fd_sc_hd__xor2_4 _29089_ (.A(_12398_),
    .B(_12403_),
    .X(_12404_));
 sky130_fd_sc_hd__xor2_4 _29090_ (.A(_12396_),
    .B(_12404_),
    .X(_12405_));
 sky130_fd_sc_hd__xnor2_4 _29091_ (.A(_12392_),
    .B(_12405_),
    .Y(_12406_));
 sky130_fd_sc_hd__xor2_4 _29092_ (.A(_12390_),
    .B(_12406_),
    .X(_12407_));
 sky130_fd_sc_hd__xnor2_4 _29093_ (.A(_12387_),
    .B(_12407_),
    .Y(_12408_));
 sky130_fd_sc_hd__xor2_4 _29094_ (.A(_12385_),
    .B(_12408_),
    .X(_12409_));
 sky130_fd_sc_hd__xnor2_4 _29095_ (.A(_12379_),
    .B(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__xor2_4 _29096_ (.A(_12377_),
    .B(_12410_),
    .X(_12411_));
 sky130_fd_sc_hd__nor2_1 _29097_ (.A(_12301_),
    .B(_12335_),
    .Y(_12412_));
 sky130_fd_sc_hd__a21o_2 _29098_ (.A1(_12334_),
    .A2(_12303_),
    .B1(_12412_),
    .X(_12413_));
 sky130_fd_sc_hd__xnor2_4 _29099_ (.A(_12411_),
    .B(_12413_),
    .Y(_12414_));
 sky130_fd_sc_hd__xor2_4 _29100_ (.A(_12373_),
    .B(_12414_),
    .X(_12415_));
 sky130_fd_sc_hd__xnor2_2 _29101_ (.A(_12369_),
    .B(_12415_),
    .Y(_12416_));
 sky130_fd_sc_hd__nor2_4 _29102_ (.A(_12368_),
    .B(_12416_),
    .Y(_12417_));
 sky130_fd_sc_hd__and2_1 _29103_ (.A(_12416_),
    .B(_12368_),
    .X(_12418_));
 sky130_fd_sc_hd__a211o_1 _29104_ (.A1(_12349_),
    .A2(_12351_),
    .B1(_12417_),
    .C1(_12418_),
    .X(_12419_));
 sky130_fd_sc_hd__o211ai_4 _29105_ (.A1(_12417_),
    .A2(_12418_),
    .B1(_12349_),
    .C1(_12351_),
    .Y(_12420_));
 sky130_fd_sc_hd__nor2_4 _29106_ (.A(_11615_),
    .B(_12345_),
    .Y(_12421_));
 sky130_fd_sc_hd__a21o_1 _29107_ (.A1(_12419_),
    .A2(_12420_),
    .B1(_12421_),
    .X(_12422_));
 sky130_fd_sc_hd__nand3_1 _29108_ (.A(_12419_),
    .B(_12421_),
    .C(_12420_),
    .Y(_12423_));
 sky130_fd_sc_hd__nand2_1 _29109_ (.A(_12357_),
    .B(_12353_),
    .Y(_12424_));
 sky130_fd_sc_hd__a21oi_1 _29110_ (.A1(_12422_),
    .A2(_12423_),
    .B1(_12424_),
    .Y(_12425_));
 sky130_fd_sc_hd__and3_1 _29111_ (.A(_12422_),
    .B(_12423_),
    .C(_12424_),
    .X(_12426_));
 sky130_fd_sc_hd__nor2_2 _29112_ (.A(_12425_),
    .B(_12426_),
    .Y(_12427_));
 sky130_fd_sc_hd__nor3b_4 _29113_ (.A(_12203_),
    .B(_12119_),
    .C_N(_12204_),
    .Y(_12428_));
 sky130_fd_sc_hd__nand3_2 _29114_ (.A(_12428_),
    .B(_12289_),
    .C(_12362_),
    .Y(_12429_));
 sky130_fd_sc_hd__nand3_1 _29115_ (.A(_12289_),
    .B(_12284_),
    .C(_12362_),
    .Y(_12430_));
 sky130_fd_sc_hd__o21ba_1 _29116_ (.A1(_12282_),
    .A2(_12360_),
    .B1_N(_12361_),
    .X(_12431_));
 sky130_fd_sc_hd__nand2_1 _29117_ (.A(_12430_),
    .B(_12431_),
    .Y(_12432_));
 sky130_fd_sc_hd__o21bai_4 _29118_ (.A1(_12429_),
    .A2(_12129_),
    .B1_N(_12432_),
    .Y(_12433_));
 sky130_fd_sc_hd__xor2_1 _29119_ (.A(_12427_),
    .B(_12433_),
    .X(_02679_));
 sky130_fd_sc_hd__a21boi_4 _29120_ (.A1(_12420_),
    .A2(_12421_),
    .B1_N(_12419_),
    .Y(_12434_));
 sky130_fd_sc_hd__and2_1 _29121_ (.A(_12413_),
    .B(_12411_),
    .X(_12435_));
 sky130_fd_sc_hd__o21bai_1 _29122_ (.A1(_12373_),
    .A2(_12414_),
    .B1_N(_12435_),
    .Y(_12436_));
 sky130_fd_sc_hd__and2_1 _29123_ (.A(_12375_),
    .B(_12002_),
    .X(_12437_));
 sky130_fd_sc_hd__o21bai_4 _29124_ (.A1(_12033_),
    .A2(_12376_),
    .B1_N(_12437_),
    .Y(_12438_));
 sky130_fd_sc_hd__xnor2_4 _29125_ (.A(_12130_),
    .B(_12438_),
    .Y(_12439_));
 sky130_fd_sc_hd__xor2_4 _29126_ (.A(net410),
    .B(_12439_),
    .X(_12440_));
 sky130_fd_sc_hd__and2_1 _29127_ (.A(_12409_),
    .B(_12379_),
    .X(_12441_));
 sky130_fd_sc_hd__o21bai_4 _29128_ (.A1(_12377_),
    .A2(_12410_),
    .B1_N(_12441_),
    .Y(_12442_));
 sky130_fd_sc_hd__and2_1 _29129_ (.A(_12383_),
    .B(_12213_),
    .X(_12443_));
 sky130_fd_sc_hd__o21bai_4 _29130_ (.A1(_12212_),
    .A2(_12384_),
    .B1_N(_12443_),
    .Y(_12444_));
 sky130_fd_sc_hd__xor2_4 _29131_ (.A(net411),
    .B(_12444_),
    .X(_12445_));
 sky130_fd_sc_hd__xor2_4 _29132_ (.A(net412),
    .B(_12445_),
    .X(_12446_));
 sky130_fd_sc_hd__and2_1 _29133_ (.A(_12407_),
    .B(_12387_),
    .X(_12447_));
 sky130_fd_sc_hd__o21bai_4 _29134_ (.A1(_12385_),
    .A2(_12408_),
    .B1_N(_12447_),
    .Y(_12448_));
 sky130_fd_sc_hd__and2_1 _29135_ (.A(_12381_),
    .B(_12388_),
    .X(_12449_));
 sky130_fd_sc_hd__o21bai_4 _29136_ (.A1(_12380_),
    .A2(_12389_),
    .B1_N(_12449_),
    .Y(_12450_));
 sky130_fd_sc_hd__xor2_4 _29137_ (.A(_12051_),
    .B(_12450_),
    .X(_12451_));
 sky130_fd_sc_hd__xor2_4 _29138_ (.A(_12144_),
    .B(_12451_),
    .X(_12452_));
 sky130_fd_sc_hd__and2_1 _29139_ (.A(_12405_),
    .B(_12392_),
    .X(_12453_));
 sky130_fd_sc_hd__o21bai_4 _29140_ (.A1(_12390_),
    .A2(_12406_),
    .B1_N(_12453_),
    .Y(_12454_));
 sky130_fd_sc_hd__nand3b_2 _29141_ (.A_N(_12394_),
    .B(_13974_),
    .C(_08589_),
    .Y(_12455_));
 sky130_fd_sc_hd__o31ai_4 _29142_ (.A1(_12782_),
    .A2(_13982_),
    .A3(_12395_),
    .B1(_12455_),
    .Y(_12456_));
 sky130_fd_sc_hd__xnor2_4 _29143_ (.A(_12456_),
    .B(_12381_),
    .Y(_12457_));
 sky130_fd_sc_hd__xnor2_4 _29144_ (.A(_12380_),
    .B(_12457_),
    .Y(_12458_));
 sky130_fd_sc_hd__or2b_1 _29145_ (.A(_12403_),
    .B_N(_12398_),
    .X(_12459_));
 sky130_fd_sc_hd__o21ai_4 _29146_ (.A1(_12396_),
    .A2(_12404_),
    .B1(_12459_),
    .Y(_12460_));
 sky130_fd_sc_hd__nand2_4 _29147_ (.A(_12780_),
    .B(_12070_),
    .Y(_12461_));
 sky130_fd_sc_hd__xnor2_4 _29148_ (.A(_12394_),
    .B(_12461_),
    .Y(_12462_));
 sky130_fd_sc_hd__xor2_4 _29149_ (.A(_12317_),
    .B(_12462_),
    .X(_12463_));
 sky130_fd_sc_hd__nand3b_2 _29150_ (.A_N(_12400_),
    .B(_08529_),
    .C(_14294_),
    .Y(_12464_));
 sky130_fd_sc_hd__o31ai_4 _29151_ (.A1(_13969_),
    .A2(_14281_),
    .A3(_12402_),
    .B1(_12464_),
    .Y(_12465_));
 sky130_fd_sc_hd__and2_2 _29152_ (.A(_08244_),
    .B(_08588_),
    .X(_12466_));
 sky130_fd_sc_hd__nand2_2 _29153_ (.A(_13963_),
    .B(_11138_),
    .Y(_12467_));
 sky130_fd_sc_hd__and2b_1 _29154_ (.A_N(_08489_),
    .B(_08527_),
    .X(_12468_));
 sky130_fd_sc_hd__xor2_4 _29155_ (.A(_12467_),
    .B(_12468_),
    .X(_12469_));
 sky130_fd_sc_hd__xor2_4 _29156_ (.A(_12466_),
    .B(_12469_),
    .X(_12470_));
 sky130_fd_sc_hd__xor2_4 _29157_ (.A(_12465_),
    .B(_12470_),
    .X(_12471_));
 sky130_fd_sc_hd__xor2_4 _29158_ (.A(_12463_),
    .B(_12471_),
    .X(_12472_));
 sky130_fd_sc_hd__xnor2_4 _29159_ (.A(_12460_),
    .B(_12472_),
    .Y(_12473_));
 sky130_fd_sc_hd__xor2_4 _29160_ (.A(_12458_),
    .B(_12473_),
    .X(_12474_));
 sky130_fd_sc_hd__xnor2_4 _29161_ (.A(_12454_),
    .B(_12474_),
    .Y(_12475_));
 sky130_fd_sc_hd__xor2_4 _29162_ (.A(_12452_),
    .B(_12475_),
    .X(_12476_));
 sky130_fd_sc_hd__xnor2_4 _29163_ (.A(_12448_),
    .B(_12476_),
    .Y(_12477_));
 sky130_fd_sc_hd__xor2_4 _29164_ (.A(_12446_),
    .B(_12477_),
    .X(_12478_));
 sky130_fd_sc_hd__xnor2_4 _29165_ (.A(_12442_),
    .B(_12478_),
    .Y(_12479_));
 sky130_fd_sc_hd__xor2_2 _29166_ (.A(_12440_),
    .B(_12479_),
    .X(_12480_));
 sky130_fd_sc_hd__or2_1 _29167_ (.A(_12436_),
    .B(_12480_),
    .X(_12481_));
 sky130_fd_sc_hd__nand2_2 _29168_ (.A(_12480_),
    .B(_12436_),
    .Y(_12482_));
 sky130_fd_sc_hd__nor2_1 _29169_ (.A(_11489_),
    .B(_12371_),
    .Y(_12483_));
 sky130_fd_sc_hd__o21ba_2 _29170_ (.A1(_12101_),
    .A2(_12372_),
    .B1_N(_12483_),
    .X(_12484_));
 sky130_fd_sc_hd__xor2_2 _29171_ (.A(_10812_),
    .B(_12484_),
    .X(_12485_));
 sky130_fd_sc_hd__and3_1 _29172_ (.A(_12481_),
    .B(_12482_),
    .C(_12485_),
    .X(_12486_));
 sky130_fd_sc_hd__a21oi_2 _29173_ (.A1(_12481_),
    .A2(_12482_),
    .B1(_12485_),
    .Y(_12487_));
 sky130_fd_sc_hd__a21o_1 _29174_ (.A1(_12415_),
    .A2(_12369_),
    .B1(_12417_),
    .X(_12488_));
 sky130_fd_sc_hd__o21bai_2 _29175_ (.A1(_12486_),
    .A2(_12487_),
    .B1_N(_12488_),
    .Y(_12489_));
 sky130_vsdinv _29176_ (.A(_12486_),
    .Y(_12490_));
 sky130_fd_sc_hd__nand3b_4 _29177_ (.A_N(_12487_),
    .B(_12488_),
    .C(_12490_),
    .Y(_12491_));
 sky130_fd_sc_hd__nor2_4 _29178_ (.A(_11615_),
    .B(_12366_),
    .Y(_12492_));
 sky130_fd_sc_hd__a21oi_4 _29179_ (.A1(_12489_),
    .A2(_12491_),
    .B1(_12492_),
    .Y(_12493_));
 sky130_fd_sc_hd__nand3_1 _29180_ (.A(_12489_),
    .B(_12491_),
    .C(_12492_),
    .Y(_12494_));
 sky130_vsdinv _29181_ (.A(_12494_),
    .Y(_12495_));
 sky130_fd_sc_hd__nor3_4 _29182_ (.A(_12434_),
    .B(_12493_),
    .C(_12495_),
    .Y(_12496_));
 sky130_fd_sc_hd__o21a_1 _29183_ (.A1(_12493_),
    .A2(_12495_),
    .B1(_12434_),
    .X(_12497_));
 sky130_fd_sc_hd__or2_1 _29184_ (.A(_12496_),
    .B(_12497_),
    .X(_12498_));
 sky130_fd_sc_hd__a21oi_1 _29185_ (.A1(_12433_),
    .A2(_12427_),
    .B1(_12426_),
    .Y(_12499_));
 sky130_fd_sc_hd__xor2_1 _29186_ (.A(_12498_),
    .B(_12499_),
    .X(_02680_));
 sky130_fd_sc_hd__a21boi_1 _29187_ (.A1(_12489_),
    .A2(_12492_),
    .B1_N(_12491_),
    .Y(_12500_));
 sky130_fd_sc_hd__and2_1 _29188_ (.A(_12438_),
    .B(_12130_),
    .X(_12501_));
 sky130_fd_sc_hd__o21bai_4 _29189_ (.A1(_12101_),
    .A2(_12439_),
    .B1_N(_12501_),
    .Y(_12502_));
 sky130_fd_sc_hd__xor2_4 _29190_ (.A(_11242_),
    .B(_12502_),
    .X(_12503_));
 sky130_fd_sc_hd__and2_1 _29191_ (.A(_12478_),
    .B(_12442_),
    .X(_12504_));
 sky130_fd_sc_hd__o21bai_4 _29192_ (.A1(_12440_),
    .A2(_12479_),
    .B1_N(_12504_),
    .Y(_12505_));
 sky130_fd_sc_hd__and2_1 _29193_ (.A(_12444_),
    .B(_12002_),
    .X(_12506_));
 sky130_fd_sc_hd__o21bai_4 _29194_ (.A1(_12033_),
    .A2(_12445_),
    .B1_N(_12506_),
    .Y(_12507_));
 sky130_fd_sc_hd__xnor2_4 _29195_ (.A(_12130_),
    .B(_12507_),
    .Y(_12508_));
 sky130_fd_sc_hd__xor2_4 _29196_ (.A(net410),
    .B(_12508_),
    .X(_12509_));
 sky130_fd_sc_hd__and2_1 _29197_ (.A(_12476_),
    .B(_12448_),
    .X(_12510_));
 sky130_fd_sc_hd__o21bai_4 _29198_ (.A1(_12446_),
    .A2(_12477_),
    .B1_N(_12510_),
    .Y(_12511_));
 sky130_fd_sc_hd__nand2_1 _29199_ (.A(_12450_),
    .B(_12213_),
    .Y(_12512_));
 sky130_fd_sc_hd__o21a_1 _29200_ (.A1(_12212_),
    .A2(_12451_),
    .B1(_12512_),
    .X(_12513_));
 sky130_fd_sc_hd__nor2_4 _29201_ (.A(_11887_),
    .B(_12513_),
    .Y(_12514_));
 sky130_fd_sc_hd__o211a_1 _29202_ (.A1(_12212_),
    .A2(_12451_),
    .B1(_11887_),
    .C1(_12512_),
    .X(_12515_));
 sky130_fd_sc_hd__a21oi_2 _29203_ (.A1(_12513_),
    .A2(_11889_),
    .B1(_11330_),
    .Y(_12516_));
 sky130_fd_sc_hd__o211ai_2 _29204_ (.A1(_12515_),
    .A2(_12514_),
    .B1(_11187_),
    .C1(_11890_),
    .Y(_12517_));
 sky130_fd_sc_hd__o31a_4 _29205_ (.A1(_12514_),
    .A2(_12515_),
    .A3(_12516_),
    .B1(_12517_),
    .X(_12518_));
 sky130_fd_sc_hd__and2_1 _29206_ (.A(_12474_),
    .B(_12454_),
    .X(_12519_));
 sky130_fd_sc_hd__o21bai_4 _29207_ (.A1(_12452_),
    .A2(_12475_),
    .B1_N(_12519_),
    .Y(_12520_));
 sky130_fd_sc_hd__nand2_1 _29208_ (.A(_12381_),
    .B(_12456_),
    .Y(_12521_));
 sky130_fd_sc_hd__o21a_2 _29209_ (.A1(_12380_),
    .A2(_12457_),
    .B1(_12521_),
    .X(_12522_));
 sky130_fd_sc_hd__xor2_4 _29210_ (.A(_12213_),
    .B(_12522_),
    .X(_12523_));
 sky130_fd_sc_hd__xor2_4 _29211_ (.A(_12144_),
    .B(_12523_),
    .X(_12524_));
 sky130_fd_sc_hd__and2_1 _29212_ (.A(_12472_),
    .B(_12460_),
    .X(_12525_));
 sky130_fd_sc_hd__o21bai_4 _29213_ (.A1(_12458_),
    .A2(_12473_),
    .B1_N(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__nand3b_2 _29214_ (.A_N(_12462_),
    .B(_12781_),
    .C(_07360_),
    .Y(_12527_));
 sky130_fd_sc_hd__o21ai_4 _29215_ (.A1(_12394_),
    .A2(_12461_),
    .B1(_12527_),
    .Y(_12528_));
 sky130_fd_sc_hd__xnor2_4 _29216_ (.A(_12231_),
    .B(_12528_),
    .Y(_12529_));
 sky130_fd_sc_hd__xnor2_4 _29217_ (.A(_12310_),
    .B(_12529_),
    .Y(_12530_));
 sky130_fd_sc_hd__or2b_1 _29218_ (.A(_12470_),
    .B_N(_12465_),
    .X(_12531_));
 sky130_fd_sc_hd__o21ai_4 _29219_ (.A1(_12463_),
    .A2(_12471_),
    .B1(_12531_),
    .Y(_12532_));
 sky130_fd_sc_hd__nand3b_2 _29220_ (.A_N(_12467_),
    .B(_08529_),
    .C(_14287_),
    .Y(_12533_));
 sky130_fd_sc_hd__o31ai_4 _29221_ (.A1(_13969_),
    .A2(_14276_),
    .A3(_12469_),
    .B1(_12533_),
    .Y(_12534_));
 sky130_fd_sc_hd__nand2_4 _29222_ (.A(_12780_),
    .B(_08244_),
    .Y(_12535_));
 sky130_fd_sc_hd__nand2_4 _29223_ (.A(_13963_),
    .B(_08596_),
    .Y(_12536_));
 sky130_fd_sc_hd__and2b_1 _29224_ (.A_N(_11138_),
    .B(_08527_),
    .X(_12537_));
 sky130_fd_sc_hd__xor2_4 _29225_ (.A(_12536_),
    .B(_12537_),
    .X(_12538_));
 sky130_fd_sc_hd__xnor2_4 _29226_ (.A(_12535_),
    .B(_12538_),
    .Y(_12539_));
 sky130_fd_sc_hd__xor2_4 _29227_ (.A(_12534_),
    .B(_12539_),
    .X(_12540_));
 sky130_fd_sc_hd__xor2_4 _29228_ (.A(_12463_),
    .B(_12540_),
    .X(_12541_));
 sky130_fd_sc_hd__xnor2_4 _29229_ (.A(_12532_),
    .B(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__xor2_4 _29230_ (.A(_12530_),
    .B(_12542_),
    .X(_12543_));
 sky130_fd_sc_hd__xnor2_4 _29231_ (.A(_12526_),
    .B(_12543_),
    .Y(_12544_));
 sky130_fd_sc_hd__xor2_4 _29232_ (.A(_12524_),
    .B(_12544_),
    .X(_12545_));
 sky130_fd_sc_hd__xnor2_4 _29233_ (.A(_12520_),
    .B(_12545_),
    .Y(_12546_));
 sky130_fd_sc_hd__xor2_4 _29234_ (.A(_12518_),
    .B(_12546_),
    .X(_12547_));
 sky130_fd_sc_hd__xnor2_4 _29235_ (.A(_12511_),
    .B(_12547_),
    .Y(_12548_));
 sky130_fd_sc_hd__xor2_4 _29236_ (.A(_12509_),
    .B(_12548_),
    .X(_12549_));
 sky130_fd_sc_hd__xor2_4 _29237_ (.A(_12505_),
    .B(_12549_),
    .X(_12550_));
 sky130_fd_sc_hd__xnor2_2 _29238_ (.A(_12503_),
    .B(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__nand3b_4 _29239_ (.A_N(_12551_),
    .B(_12482_),
    .C(_12490_),
    .Y(_12552_));
 sky130_fd_sc_hd__nor2_2 _29240_ (.A(_11615_),
    .B(_12484_),
    .Y(_12553_));
 sky130_fd_sc_hd__a21boi_1 _29241_ (.A1(_12481_),
    .A2(_12485_),
    .B1_N(_12482_),
    .Y(_12554_));
 sky130_vsdinv _29242_ (.A(_12554_),
    .Y(_12555_));
 sky130_fd_sc_hd__nand2_4 _29243_ (.A(_12551_),
    .B(_12555_),
    .Y(_12556_));
 sky130_fd_sc_hd__nand3_4 _29244_ (.A(_12552_),
    .B(_12553_),
    .C(_12556_),
    .Y(_12557_));
 sky130_fd_sc_hd__o2bb2ai_1 _29245_ (.A1_N(_12556_),
    .A2_N(_12552_),
    .B1(_11615_),
    .B2(_12484_),
    .Y(_12558_));
 sky130_fd_sc_hd__and3b_1 _29246_ (.A_N(_12500_),
    .B(_12557_),
    .C(_12558_),
    .X(_12559_));
 sky130_vsdinv _29247_ (.A(_12559_),
    .Y(_12560_));
 sky130_fd_sc_hd__a21bo_1 _29248_ (.A1(_12558_),
    .A2(_12557_),
    .B1_N(_12500_),
    .X(_12561_));
 sky130_fd_sc_hd__nand2_4 _29249_ (.A(_12560_),
    .B(_12561_),
    .Y(_12562_));
 sky130_fd_sc_hd__nor3b_4 _29250_ (.A(_12496_),
    .B(_12497_),
    .C_N(_12427_),
    .Y(_12563_));
 sky130_fd_sc_hd__o21ba_1 _29251_ (.A1(_12426_),
    .A2(_12496_),
    .B1_N(_12497_),
    .X(_12564_));
 sky130_fd_sc_hd__a21oi_4 _29252_ (.A1(_12433_),
    .A2(_12563_),
    .B1(_12564_),
    .Y(_12565_));
 sky130_fd_sc_hd__xor2_4 _29253_ (.A(_12562_),
    .B(_12565_),
    .X(_02681_));
 sky130_fd_sc_hd__o21bai_1 _29254_ (.A1(_12562_),
    .A2(_12565_),
    .B1_N(_12559_),
    .Y(_12566_));
 sky130_fd_sc_hd__and2_1 _29255_ (.A(_12541_),
    .B(_12532_),
    .X(_12567_));
 sky130_fd_sc_hd__o21bai_1 _29256_ (.A1(_12530_),
    .A2(_12542_),
    .B1_N(_12567_),
    .Y(_12568_));
 sky130_fd_sc_hd__and2_1 _29257_ (.A(_12545_),
    .B(_12520_),
    .X(_12569_));
 sky130_fd_sc_hd__o21bai_1 _29258_ (.A1(_12518_),
    .A2(_12546_),
    .B1_N(_12569_),
    .Y(_12570_));
 sky130_fd_sc_hd__xor2_1 _29259_ (.A(_12568_),
    .B(_12570_),
    .X(_12571_));
 sky130_fd_sc_hd__xnor2_1 _29260_ (.A(_12535_),
    .B(_12571_),
    .Y(_12572_));
 sky130_fd_sc_hd__and2_1 _29261_ (.A(_12781_),
    .B(_13963_),
    .X(_12573_));
 sky130_vsdinv _29262_ (.A(_12573_),
    .Y(_12574_));
 sky130_fd_sc_hd__or2b_1 _29263_ (.A(_12539_),
    .B_N(_12534_),
    .X(_12575_));
 sky130_fd_sc_hd__o21a_1 _29264_ (.A1(_12463_),
    .A2(_12540_),
    .B1(_12575_),
    .X(_12576_));
 sky130_fd_sc_hd__and2b_1 _29265_ (.A_N(_12503_),
    .B(_12550_),
    .X(_12577_));
 sky130_fd_sc_hd__a211o_1 _29266_ (.A1(_12549_),
    .A2(_12505_),
    .B1(_12576_),
    .C1(_12577_),
    .X(_12578_));
 sky130_fd_sc_hd__and2_1 _29267_ (.A(_12549_),
    .B(_12505_),
    .X(_12579_));
 sky130_fd_sc_hd__o21ai_2 _29268_ (.A1(_12579_),
    .A2(_12577_),
    .B1(_12576_),
    .Y(_12580_));
 sky130_fd_sc_hd__nor2_2 _29269_ (.A(_12514_),
    .B(_12516_),
    .Y(_12581_));
 sky130_fd_sc_hd__mux2_2 _29270_ (.A0(_11356_),
    .A1(_11358_),
    .S(_09978_),
    .X(_12582_));
 sky130_fd_sc_hd__xor2_2 _29271_ (.A(_12581_),
    .B(_12582_),
    .X(_12583_));
 sky130_vsdinv _29272_ (.A(_12583_),
    .Y(_12584_));
 sky130_fd_sc_hd__a21oi_4 _29273_ (.A1(_12578_),
    .A2(_12580_),
    .B1(_12584_),
    .Y(_12585_));
 sky130_fd_sc_hd__and3_1 _29274_ (.A(_12578_),
    .B(_12580_),
    .C(_12584_),
    .X(_12586_));
 sky130_fd_sc_hd__nor3_4 _29275_ (.A(_12574_),
    .B(_12585_),
    .C(_12586_),
    .Y(_12587_));
 sky130_fd_sc_hd__o21a_1 _29276_ (.A1(_12585_),
    .A2(_12586_),
    .B1(_12574_),
    .X(_12588_));
 sky130_fd_sc_hd__nor3_2 _29277_ (.A(_12572_),
    .B(_12587_),
    .C(_12588_),
    .Y(_12589_));
 sky130_fd_sc_hd__o21a_1 _29278_ (.A1(_12587_),
    .A2(_12588_),
    .B1(_12572_),
    .X(_12590_));
 sky130_fd_sc_hd__or2_1 _29279_ (.A(_12589_),
    .B(_12590_),
    .X(_12591_));
 sky130_fd_sc_hd__nand2_1 _29280_ (.A(_12543_),
    .B(_12526_),
    .Y(_12592_));
 sky130_fd_sc_hd__o21a_1 _29281_ (.A1(_12524_),
    .A2(_12544_),
    .B1(_12592_),
    .X(_12593_));
 sky130_fd_sc_hd__a21bo_1 _29282_ (.A1(_12557_),
    .A2(_12556_),
    .B1_N(_12593_),
    .X(_12594_));
 sky130_fd_sc_hd__nand3b_2 _29283_ (.A_N(_12593_),
    .B(_12557_),
    .C(_12556_),
    .Y(_12595_));
 sky130_fd_sc_hd__o21a_1 _29284_ (.A1(_12047_),
    .A2(_12522_),
    .B1(_11840_),
    .X(_12596_));
 sky130_fd_sc_hd__a21o_1 _29285_ (.A1(_12142_),
    .A2(_12522_),
    .B1(_12596_),
    .X(_12597_));
 sky130_fd_sc_hd__a21o_1 _29286_ (.A1(_12594_),
    .A2(_12595_),
    .B1(_12597_),
    .X(_12598_));
 sky130_fd_sc_hd__nand3_2 _29287_ (.A(_12594_),
    .B(_12597_),
    .C(_12595_),
    .Y(_12599_));
 sky130_fd_sc_hd__and2_2 _29288_ (.A(_12529_),
    .B(_12380_),
    .X(_12600_));
 sky130_fd_sc_hd__nand2_2 _29289_ (.A(_14277_),
    .B(_08529_),
    .Y(_12601_));
 sky130_fd_sc_hd__nand2_1 _29290_ (.A(_12507_),
    .B(_12130_),
    .Y(_12602_));
 sky130_fd_sc_hd__o21a_2 _29291_ (.A1(_12101_),
    .A2(_12508_),
    .B1(_12602_),
    .X(_12603_));
 sky130_fd_sc_hd__nor3_2 _29292_ (.A(_08482_),
    .B(_12806_),
    .C(_12536_),
    .Y(_12604_));
 sky130_fd_sc_hd__o21ba_2 _29293_ (.A1(_12535_),
    .A2(_12538_),
    .B1_N(_12604_),
    .X(_12605_));
 sky130_fd_sc_hd__nor2_4 _29294_ (.A(_10813_),
    .B(_12502_),
    .Y(_12606_));
 sky130_fd_sc_hd__xor2_4 _29295_ (.A(_12605_),
    .B(_12606_),
    .X(_12607_));
 sky130_fd_sc_hd__xor2_4 _29296_ (.A(_12603_),
    .B(_12607_),
    .X(_12608_));
 sky130_fd_sc_hd__xor2_4 _29297_ (.A(_12601_),
    .B(_12608_),
    .X(_12609_));
 sky130_fd_sc_hd__xor2_4 _29298_ (.A(_12600_),
    .B(_12609_),
    .X(_12610_));
 sky130_fd_sc_hd__and2_2 _29299_ (.A(_12528_),
    .B(_12381_),
    .X(_12611_));
 sky130_fd_sc_hd__and2_1 _29300_ (.A(_12547_),
    .B(_12511_),
    .X(_12612_));
 sky130_fd_sc_hd__o21bai_4 _29301_ (.A1(_12509_),
    .A2(_12548_),
    .B1_N(_12612_),
    .Y(_12613_));
 sky130_fd_sc_hd__xor2_4 _29302_ (.A(_12463_),
    .B(_12613_),
    .X(_12614_));
 sky130_fd_sc_hd__xor2_4 _29303_ (.A(_12611_),
    .B(_12614_),
    .X(_12615_));
 sky130_fd_sc_hd__xor2_4 _29304_ (.A(_12610_),
    .B(_12615_),
    .X(_12616_));
 sky130_fd_sc_hd__a21o_1 _29305_ (.A1(_12598_),
    .A2(_12599_),
    .B1(_12616_),
    .X(_12617_));
 sky130_fd_sc_hd__nand3_2 _29306_ (.A(_12598_),
    .B(_12616_),
    .C(_12599_),
    .Y(_12618_));
 sky130_fd_sc_hd__nand2_1 _29307_ (.A(_12617_),
    .B(_12618_),
    .Y(_12619_));
 sky130_fd_sc_hd__xor2_1 _29308_ (.A(_12591_),
    .B(_12619_),
    .X(_12620_));
 sky130_fd_sc_hd__nand2_2 _29309_ (.A(_12566_),
    .B(_12620_),
    .Y(_12621_));
 sky130_fd_sc_hd__a21oi_1 _29310_ (.A1(_12617_),
    .A2(_12618_),
    .B1(_12591_),
    .Y(_12622_));
 sky130_fd_sc_hd__o211a_1 _29311_ (.A1(_12590_),
    .A2(_12589_),
    .B1(_12618_),
    .C1(_12617_),
    .X(_12623_));
 sky130_fd_sc_hd__nor2_2 _29312_ (.A(_12622_),
    .B(_12623_),
    .Y(_12624_));
 sky130_fd_sc_hd__o211ai_4 _29313_ (.A1(_12562_),
    .A2(_12565_),
    .B1(_12560_),
    .C1(_12624_),
    .Y(_12625_));
 sky130_fd_sc_hd__nand2_8 _29314_ (.A(_12621_),
    .B(_12625_),
    .Y(_02682_));
 sky130_fd_sc_hd__a21oi_1 _29315_ (.A1(_04945_),
    .A2(_04919_),
    .B1(_05020_),
    .Y(_12626_));
 sky130_fd_sc_hd__xor2_1 _29316_ (.A(_05025_),
    .B(_12626_),
    .X(_02628_));
 sky130_fd_sc_hd__and2_1 _29317_ (.A(_00049_),
    .B(_02321_),
    .X(_00050_));
 sky130_fd_sc_hd__nor3b_1 _29318_ (.A(_14646_),
    .B(_13838_),
    .C_N(_00066_),
    .Y(_00068_));
 sky130_fd_sc_hd__nor2b_1 _29319_ (.A(_14646_),
    .B_N(_00084_),
    .Y(_00085_));
 sky130_fd_sc_hd__nor2b_1 _29320_ (.A(_14646_),
    .B_N(_00094_),
    .Y(_00095_));
 sky130_fd_sc_hd__o21a_4 _29321_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(_12797_),
    .X(_00216_));
 sky130_fd_sc_hd__a21boi_2 _29322_ (.A1(_04398_),
    .A2(_12866_),
    .B1_N(_00321_),
    .Y(_12627_));
 sky130_fd_sc_hd__o211ai_2 _29323_ (.A1(_12878_),
    .A2(_13101_),
    .B1(_12917_),
    .C1(_00321_),
    .Y(_12628_));
 sky130_fd_sc_hd__o211a_1 _29324_ (.A1(_14651_),
    .A2(_12627_),
    .B1(_13542_),
    .C1(_12628_),
    .X(_04072_));
 sky130_fd_sc_hd__conb_1 _29325_ (.LO(net134));
 sky130_fd_sc_hd__conb_1 _29326_ (.LO(net145));
 sky130_fd_sc_hd__conb_1 _29327_ (.LO(net167));
 sky130_fd_sc_hd__conb_1 _29328_ (.LO(net178));
 sky130_fd_sc_hd__conb_1 _29329_ (.LO(net371));
 sky130_fd_sc_hd__conb_1 _29330_ (.LO(net382));
 sky130_fd_sc_hd__conb_1 _29331_ (.LO(net393));
 sky130_fd_sc_hd__conb_1 _29332_ (.LO(net400));
 sky130_fd_sc_hd__conb_1 _29333_ (.LO(net401));
 sky130_fd_sc_hd__conb_1 _29334_ (.LO(net402));
 sky130_fd_sc_hd__conb_1 _29335_ (.LO(net403));
 sky130_fd_sc_hd__conb_1 _29336_ (.LO(net404));
 sky130_fd_sc_hd__conb_1 _29337_ (.LO(net405));
 sky130_fd_sc_hd__conb_1 _29338_ (.LO(net406));
 sky130_fd_sc_hd__conb_1 _29339_ (.LO(net372));
 sky130_fd_sc_hd__conb_1 _29340_ (.LO(net373));
 sky130_fd_sc_hd__conb_1 _29341_ (.LO(net374));
 sky130_fd_sc_hd__conb_1 _29342_ (.LO(net375));
 sky130_fd_sc_hd__conb_1 _29343_ (.LO(net376));
 sky130_fd_sc_hd__conb_1 _29344_ (.LO(net377));
 sky130_fd_sc_hd__conb_1 _29345_ (.LO(net378));
 sky130_fd_sc_hd__conb_1 _29346_ (.LO(net379));
 sky130_fd_sc_hd__conb_1 _29347_ (.LO(net380));
 sky130_fd_sc_hd__conb_1 _29348_ (.LO(net381));
 sky130_fd_sc_hd__conb_1 _29349_ (.LO(net383));
 sky130_fd_sc_hd__conb_1 _29350_ (.LO(net384));
 sky130_fd_sc_hd__conb_1 _29351_ (.LO(net385));
 sky130_fd_sc_hd__conb_1 _29352_ (.LO(net386));
 sky130_fd_sc_hd__conb_1 _29353_ (.LO(net387));
 sky130_fd_sc_hd__conb_1 _29354_ (.LO(net388));
 sky130_fd_sc_hd__conb_1 _29355_ (.LO(net389));
 sky130_fd_sc_hd__conb_1 _29356_ (.LO(net390));
 sky130_fd_sc_hd__conb_1 _29357_ (.LO(net391));
 sky130_fd_sc_hd__conb_1 _29358_ (.LO(net392));
 sky130_fd_sc_hd__conb_1 _29359_ (.LO(net394));
 sky130_fd_sc_hd__conb_1 _29360_ (.LO(net395));
 sky130_fd_sc_hd__conb_1 _29361_ (.LO(net396));
 sky130_fd_sc_hd__conb_1 _29362_ (.LO(net397));
 sky130_fd_sc_hd__conb_1 _29363_ (.LO(net398));
 sky130_fd_sc_hd__conb_1 _29364_ (.LO(net399));
 sky130_fd_sc_hd__conb_1 _29365_ (.LO(net407));
 sky130_fd_sc_hd__conb_1 _29366_ (.LO(_00313_));
 sky130_fd_sc_hd__clkbuf_4 _29367_ (.A(net200),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 _29368_ (.A(net211),
    .X(net349));
 sky130_fd_sc_hd__buf_4 _29369_ (.A(net490),
    .X(net360));
 sky130_fd_sc_hd__buf_2 _29370_ (.A(net489),
    .X(net363));
 sky130_fd_sc_hd__buf_4 _29371_ (.A(net226),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 _29372_ (.A(net227),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 _29373_ (.A(net228),
    .X(net366));
 sky130_fd_sc_hd__buf_1 _29374_ (.A(net229),
    .X(net367));
 sky130_fd_sc_hd__mux2_8 _29375_ (.A0(decoder_trigger),
    .A1(_02410_),
    .S(_00309_),
    .X(_15209_));
 sky130_fd_sc_hd__mux2_1 _29376_ (.A0(\reg_out[2] ),
    .A1(\reg_next_pc[2] ),
    .S(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_8 _29377_ (.A0(_02184_),
    .A1(net328),
    .S(net442),
    .X(net189));
 sky130_fd_sc_hd__mux2_1 _29378_ (.A0(\reg_out[3] ),
    .A1(\reg_next_pc[3] ),
    .S(_02183_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_4 _29379_ (.A0(_02185_),
    .A1(net331),
    .S(net441),
    .X(net192));
 sky130_fd_sc_hd__mux2_1 _29380_ (.A0(\reg_out[4] ),
    .A1(\reg_next_pc[4] ),
    .S(_02183_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_8 _29381_ (.A0(_02186_),
    .A1(net332),
    .S(net443),
    .X(net193));
 sky130_fd_sc_hd__mux2_1 _29382_ (.A0(\reg_out[5] ),
    .A1(\reg_next_pc[5] ),
    .S(_02183_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_8 _29383_ (.A0(_02187_),
    .A1(net333),
    .S(net443),
    .X(net194));
 sky130_fd_sc_hd__mux2_1 _29384_ (.A0(\reg_out[6] ),
    .A1(\reg_next_pc[6] ),
    .S(_02183_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_4 _29385_ (.A0(_02188_),
    .A1(net334),
    .S(net441),
    .X(net195));
 sky130_fd_sc_hd__mux2_2 _29386_ (.A0(\reg_out[7] ),
    .A1(\reg_next_pc[7] ),
    .S(_02183_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_4 _29387_ (.A0(_02189_),
    .A1(net335),
    .S(net441),
    .X(net196));
 sky130_fd_sc_hd__mux2_1 _29388_ (.A0(\reg_out[8] ),
    .A1(\reg_next_pc[8] ),
    .S(_02183_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_4 _29389_ (.A0(_02190_),
    .A1(net336),
    .S(net441),
    .X(net197));
 sky130_fd_sc_hd__mux2_1 _29390_ (.A0(\reg_out[9] ),
    .A1(\reg_next_pc[9] ),
    .S(_02183_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_8 _29391_ (.A0(_02191_),
    .A1(net337),
    .S(net442),
    .X(net198));
 sky130_fd_sc_hd__mux2_1 _29392_ (.A0(\reg_out[10] ),
    .A1(\reg_next_pc[10] ),
    .S(_02183_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_8 _29393_ (.A0(_02192_),
    .A1(net307),
    .S(net441),
    .X(net168));
 sky130_fd_sc_hd__mux2_2 _29394_ (.A0(\reg_out[11] ),
    .A1(\reg_next_pc[11] ),
    .S(_02183_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_8 _29395_ (.A0(_02193_),
    .A1(net308),
    .S(net440),
    .X(net169));
 sky130_fd_sc_hd__mux2_1 _29396_ (.A0(\reg_out[12] ),
    .A1(\reg_next_pc[12] ),
    .S(_02183_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_8 _29397_ (.A0(_02194_),
    .A1(net309),
    .S(net440),
    .X(net170));
 sky130_fd_sc_hd__mux2_2 _29398_ (.A0(\reg_out[13] ),
    .A1(\reg_next_pc[13] ),
    .S(_02183_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_8 _29399_ (.A0(_02195_),
    .A1(net310),
    .S(net441),
    .X(net171));
 sky130_fd_sc_hd__mux2_1 _29400_ (.A0(\reg_out[14] ),
    .A1(\reg_next_pc[14] ),
    .S(_02183_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_8 _29401_ (.A0(_02196_),
    .A1(net311),
    .S(net442),
    .X(net172));
 sky130_fd_sc_hd__mux2_1 _29402_ (.A0(\reg_out[15] ),
    .A1(\reg_next_pc[15] ),
    .S(_02183_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_2 _29403_ (.A0(_02197_),
    .A1(net312),
    .S(net440),
    .X(net173));
 sky130_fd_sc_hd__mux2_1 _29404_ (.A0(\reg_out[16] ),
    .A1(\reg_next_pc[16] ),
    .S(_02183_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_8 _29405_ (.A0(_02198_),
    .A1(net313),
    .S(net442),
    .X(net174));
 sky130_fd_sc_hd__mux2_2 _29406_ (.A0(\reg_out[17] ),
    .A1(\reg_next_pc[17] ),
    .S(_02183_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_8 _29407_ (.A0(_02199_),
    .A1(net314),
    .S(net443),
    .X(net175));
 sky130_fd_sc_hd__mux2_2 _29408_ (.A0(\reg_out[18] ),
    .A1(\reg_next_pc[18] ),
    .S(_02183_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_8 _29409_ (.A0(_02200_),
    .A1(net315),
    .S(net440),
    .X(net176));
 sky130_fd_sc_hd__mux2_1 _29410_ (.A0(\reg_out[19] ),
    .A1(\reg_next_pc[19] ),
    .S(_02183_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_8 _29411_ (.A0(_02201_),
    .A1(net316),
    .S(net442),
    .X(net177));
 sky130_fd_sc_hd__mux2_2 _29412_ (.A0(\reg_out[20] ),
    .A1(\reg_next_pc[20] ),
    .S(_02183_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_4 _29413_ (.A0(_02202_),
    .A1(net318),
    .S(net440),
    .X(net179));
 sky130_fd_sc_hd__mux2_2 _29414_ (.A0(\reg_out[21] ),
    .A1(\reg_next_pc[21] ),
    .S(_02183_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_8 _29415_ (.A0(_02203_),
    .A1(net319),
    .S(net443),
    .X(net180));
 sky130_fd_sc_hd__mux2_2 _29416_ (.A0(\reg_out[22] ),
    .A1(\reg_next_pc[22] ),
    .S(_02183_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_8 _29417_ (.A0(_02204_),
    .A1(net320),
    .S(net443),
    .X(net181));
 sky130_fd_sc_hd__mux2_2 _29418_ (.A0(\reg_out[23] ),
    .A1(\reg_next_pc[23] ),
    .S(_02183_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_8 _29419_ (.A0(_02205_),
    .A1(net321),
    .S(net440),
    .X(net182));
 sky130_fd_sc_hd__mux2_2 _29420_ (.A0(\reg_out[24] ),
    .A1(\reg_next_pc[24] ),
    .S(_02183_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_8 _29421_ (.A0(_02206_),
    .A1(net322),
    .S(net441),
    .X(net183));
 sky130_fd_sc_hd__mux2_2 _29422_ (.A0(\reg_out[25] ),
    .A1(\reg_next_pc[25] ),
    .S(_02183_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_4 _29423_ (.A0(_02207_),
    .A1(net323),
    .S(net440),
    .X(net184));
 sky130_fd_sc_hd__mux2_2 _29424_ (.A0(\reg_out[26] ),
    .A1(\reg_next_pc[26] ),
    .S(_02183_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_8 _29425_ (.A0(_02208_),
    .A1(net324),
    .S(net440),
    .X(net185));
 sky130_fd_sc_hd__mux2_1 _29426_ (.A0(\reg_out[27] ),
    .A1(\reg_next_pc[27] ),
    .S(_02183_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_4 _29427_ (.A0(_02209_),
    .A1(net325),
    .S(_00301_),
    .X(net186));
 sky130_fd_sc_hd__mux2_2 _29428_ (.A0(\reg_out[28] ),
    .A1(\reg_next_pc[28] ),
    .S(_02183_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_8 _29429_ (.A0(_02210_),
    .A1(net326),
    .S(net440),
    .X(net187));
 sky130_fd_sc_hd__mux2_1 _29430_ (.A0(\reg_out[29] ),
    .A1(\reg_next_pc[29] ),
    .S(_02183_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_8 _29431_ (.A0(_02211_),
    .A1(net327),
    .S(net443),
    .X(net188));
 sky130_fd_sc_hd__mux2_1 _29432_ (.A0(\reg_out[30] ),
    .A1(\reg_next_pc[30] ),
    .S(_02183_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_8 _29433_ (.A0(_02212_),
    .A1(net329),
    .S(_00301_),
    .X(net190));
 sky130_fd_sc_hd__mux2_2 _29434_ (.A0(\reg_out[31] ),
    .A1(\reg_next_pc[31] ),
    .S(_02183_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_4 _29435_ (.A0(_02213_),
    .A1(net330),
    .S(net441),
    .X(net191));
 sky130_fd_sc_hd__mux2_8 _29436_ (.A0(_02167_),
    .A1(net368),
    .S(net450),
    .X(net230));
 sky130_fd_sc_hd__mux2_8 _29437_ (.A0(_02168_),
    .A1(net369),
    .S(net450),
    .X(net231));
 sky130_fd_sc_hd__mux2_8 _29438_ (.A0(_02169_),
    .A1(net339),
    .S(net450),
    .X(net201));
 sky130_fd_sc_hd__mux2_4 _29439_ (.A0(_02170_),
    .A1(net340),
    .S(net452),
    .X(net202));
 sky130_fd_sc_hd__mux2_8 _29440_ (.A0(_02171_),
    .A1(net341),
    .S(net451),
    .X(net203));
 sky130_fd_sc_hd__mux2_8 _29441_ (.A0(_02172_),
    .A1(net342),
    .S(net452),
    .X(net204));
 sky130_fd_sc_hd__mux2_8 _29442_ (.A0(_02173_),
    .A1(net343),
    .S(net451),
    .X(net205));
 sky130_fd_sc_hd__mux2_8 _29443_ (.A0(_02174_),
    .A1(net344),
    .S(net451),
    .X(net206));
 sky130_fd_sc_hd__mux2_8 _29444_ (.A0(_02175_),
    .A1(net345),
    .S(net452),
    .X(net207));
 sky130_fd_sc_hd__mux2_8 _29445_ (.A0(_02176_),
    .A1(net346),
    .S(net451),
    .X(net208));
 sky130_fd_sc_hd__mux2_8 _29446_ (.A0(_02177_),
    .A1(net347),
    .S(net450),
    .X(net209));
 sky130_fd_sc_hd__mux2_8 _29447_ (.A0(_02178_),
    .A1(net348),
    .S(net450),
    .X(net210));
 sky130_fd_sc_hd__mux2_8 _29448_ (.A0(_02179_),
    .A1(net350),
    .S(net450),
    .X(net212));
 sky130_fd_sc_hd__mux2_4 _29449_ (.A0(_02180_),
    .A1(net351),
    .S(net451),
    .X(net213));
 sky130_fd_sc_hd__mux2_8 _29450_ (.A0(_02181_),
    .A1(net352),
    .S(net451),
    .X(net214));
 sky130_fd_sc_hd__mux2_8 _29451_ (.A0(_02182_),
    .A1(net353),
    .S(net451),
    .X(net215));
 sky130_fd_sc_hd__mux2_8 _29452_ (.A0(_02167_),
    .A1(net354),
    .S(net450),
    .X(net216));
 sky130_fd_sc_hd__mux2_8 _29453_ (.A0(_02168_),
    .A1(net355),
    .S(net450),
    .X(net217));
 sky130_fd_sc_hd__mux2_8 _29454_ (.A0(_02169_),
    .A1(net356),
    .S(net450),
    .X(net218));
 sky130_fd_sc_hd__mux2_8 _29455_ (.A0(_02170_),
    .A1(net357),
    .S(net452),
    .X(net219));
 sky130_fd_sc_hd__mux2_8 _29456_ (.A0(_02171_),
    .A1(net358),
    .S(net451),
    .X(net220));
 sky130_fd_sc_hd__mux2_4 _29457_ (.A0(_02172_),
    .A1(net359),
    .S(net452),
    .X(net221));
 sky130_fd_sc_hd__mux2_8 _29458_ (.A0(_02173_),
    .A1(net361),
    .S(net451),
    .X(net223));
 sky130_fd_sc_hd__mux2_8 _29459_ (.A0(_02174_),
    .A1(net362),
    .S(net451),
    .X(net224));
 sky130_fd_sc_hd__mux2_1 _29460_ (.A0(\mem_rdata_q[7] ),
    .A1(net62),
    .S(mem_xfer),
    .X(\mem_rdata_latched[7] ));
 sky130_fd_sc_hd__mux2_1 _29461_ (.A0(\mem_rdata_q[8] ),
    .A1(net63),
    .S(net445),
    .X(\mem_rdata_latched[8] ));
 sky130_fd_sc_hd__mux2_1 _29462_ (.A0(\mem_rdata_q[9] ),
    .A1(net64),
    .S(net445),
    .X(\mem_rdata_latched[9] ));
 sky130_fd_sc_hd__mux2_1 _29463_ (.A0(\mem_rdata_q[10] ),
    .A1(net34),
    .S(net445),
    .X(\mem_rdata_latched[10] ));
 sky130_fd_sc_hd__mux2_1 _29464_ (.A0(\mem_rdata_q[11] ),
    .A1(net35),
    .S(net444),
    .X(\mem_rdata_latched[11] ));
 sky130_fd_sc_hd__mux2_2 _29465_ (.A0(\mem_rdata_q[12] ),
    .A1(net36),
    .S(net445),
    .X(\mem_rdata_latched[12] ));
 sky130_fd_sc_hd__mux2_2 _29466_ (.A0(\mem_rdata_q[13] ),
    .A1(net37),
    .S(net445),
    .X(\mem_rdata_latched[13] ));
 sky130_fd_sc_hd__mux2_2 _29467_ (.A0(\mem_rdata_q[14] ),
    .A1(net38),
    .S(net445),
    .X(\mem_rdata_latched[14] ));
 sky130_fd_sc_hd__mux2_1 _29468_ (.A0(\mem_rdata_q[15] ),
    .A1(net500),
    .S(net444),
    .X(\mem_rdata_latched[15] ));
 sky130_fd_sc_hd__mux2_1 _29469_ (.A0(\mem_rdata_q[16] ),
    .A1(net40),
    .S(net444),
    .X(\mem_rdata_latched[16] ));
 sky130_fd_sc_hd__mux2_1 _29470_ (.A0(\mem_rdata_q[17] ),
    .A1(net499),
    .S(net444),
    .X(\mem_rdata_latched[17] ));
 sky130_fd_sc_hd__mux2_1 _29471_ (.A0(\mem_rdata_q[18] ),
    .A1(net42),
    .S(net444),
    .X(\mem_rdata_latched[18] ));
 sky130_fd_sc_hd__mux2_1 _29472_ (.A0(\mem_rdata_q[19] ),
    .A1(net498),
    .S(net444),
    .X(\mem_rdata_latched[19] ));
 sky130_fd_sc_hd__mux2_1 _29473_ (.A0(\mem_rdata_q[20] ),
    .A1(net45),
    .S(net445),
    .X(\mem_rdata_latched[20] ));
 sky130_fd_sc_hd__mux2_1 _29474_ (.A0(\mem_rdata_q[21] ),
    .A1(net46),
    .S(net444),
    .X(\mem_rdata_latched[21] ));
 sky130_fd_sc_hd__mux2_1 _29475_ (.A0(\mem_rdata_q[22] ),
    .A1(net47),
    .S(net444),
    .X(\mem_rdata_latched[22] ));
 sky130_fd_sc_hd__mux2_1 _29476_ (.A0(\mem_rdata_q[23] ),
    .A1(net48),
    .S(net444),
    .X(\mem_rdata_latched[23] ));
 sky130_fd_sc_hd__mux2_1 _29477_ (.A0(\mem_rdata_q[24] ),
    .A1(net49),
    .S(net444),
    .X(\mem_rdata_latched[24] ));
 sky130_fd_sc_hd__mux2_2 _29478_ (.A0(\mem_rdata_q[25] ),
    .A1(net50),
    .S(net444),
    .X(\mem_rdata_latched[25] ));
 sky130_fd_sc_hd__mux2_2 _29479_ (.A0(\mem_rdata_q[26] ),
    .A1(net51),
    .S(net444),
    .X(\mem_rdata_latched[26] ));
 sky130_fd_sc_hd__mux2_2 _29480_ (.A0(\mem_rdata_q[27] ),
    .A1(net52),
    .S(net444),
    .X(\mem_rdata_latched[27] ));
 sky130_fd_sc_hd__mux2_2 _29481_ (.A0(\mem_rdata_q[28] ),
    .A1(net53),
    .S(net444),
    .X(\mem_rdata_latched[28] ));
 sky130_fd_sc_hd__mux2_1 _29482_ (.A0(\mem_rdata_q[29] ),
    .A1(net54),
    .S(net445),
    .X(\mem_rdata_latched[29] ));
 sky130_fd_sc_hd__mux2_1 _29483_ (.A0(\mem_rdata_q[30] ),
    .A1(net497),
    .S(net445),
    .X(\mem_rdata_latched[30] ));
 sky130_fd_sc_hd__mux2_4 _29484_ (.A0(\mem_rdata_q[31] ),
    .A1(net57),
    .S(net445),
    .X(\mem_rdata_latched[31] ));
 sky130_fd_sc_hd__mux2_1 _29485_ (.A0(_02134_),
    .A1(\alu_add_sub[0] ),
    .S(_02133_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__mux2_1 _29486_ (.A0(_02135_),
    .A1(\alu_add_sub[1] ),
    .S(_02133_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__mux2_1 _29487_ (.A0(_02136_),
    .A1(\alu_add_sub[2] ),
    .S(_02133_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__mux2_1 _29488_ (.A0(_02137_),
    .A1(\alu_add_sub[3] ),
    .S(_02133_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__mux2_1 _29489_ (.A0(_02138_),
    .A1(\alu_add_sub[4] ),
    .S(_02133_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__mux2_1 _29490_ (.A0(_02139_),
    .A1(\alu_add_sub[5] ),
    .S(_02133_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__mux2_1 _29491_ (.A0(_02140_),
    .A1(\alu_add_sub[6] ),
    .S(_02133_),
    .X(\alu_out[6] ));
 sky130_fd_sc_hd__mux2_1 _29492_ (.A0(_02141_),
    .A1(\alu_add_sub[7] ),
    .S(_02133_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__mux2_1 _29493_ (.A0(_02142_),
    .A1(\alu_add_sub[8] ),
    .S(_02133_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__mux2_1 _29494_ (.A0(_02143_),
    .A1(\alu_add_sub[9] ),
    .S(_02133_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__mux2_1 _29495_ (.A0(_02144_),
    .A1(\alu_add_sub[10] ),
    .S(_02133_),
    .X(\alu_out[10] ));
 sky130_fd_sc_hd__mux2_1 _29496_ (.A0(_02145_),
    .A1(\alu_add_sub[11] ),
    .S(_02133_),
    .X(\alu_out[11] ));
 sky130_fd_sc_hd__mux2_2 _29497_ (.A0(_02146_),
    .A1(\alu_add_sub[12] ),
    .S(_02133_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__mux2_1 _29498_ (.A0(_02147_),
    .A1(\alu_add_sub[13] ),
    .S(_02133_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__mux2_1 _29499_ (.A0(_02148_),
    .A1(\alu_add_sub[14] ),
    .S(_02133_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__mux2_1 _29500_ (.A0(_02149_),
    .A1(\alu_add_sub[15] ),
    .S(_02133_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__mux2_1 _29501_ (.A0(_02150_),
    .A1(\alu_add_sub[16] ),
    .S(_02133_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__mux2_1 _29502_ (.A0(_02151_),
    .A1(\alu_add_sub[17] ),
    .S(_02133_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__mux2_1 _29503_ (.A0(_02152_),
    .A1(\alu_add_sub[18] ),
    .S(_02133_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__mux2_1 _29504_ (.A0(_02153_),
    .A1(\alu_add_sub[19] ),
    .S(_02133_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__mux2_2 _29505_ (.A0(_02154_),
    .A1(\alu_add_sub[20] ),
    .S(_02133_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__mux2_1 _29506_ (.A0(_02155_),
    .A1(\alu_add_sub[21] ),
    .S(_02133_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__mux2_1 _29507_ (.A0(_02156_),
    .A1(\alu_add_sub[22] ),
    .S(_02133_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__mux2_2 _29508_ (.A0(_02157_),
    .A1(\alu_add_sub[23] ),
    .S(_02133_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__mux2_2 _29509_ (.A0(_02158_),
    .A1(\alu_add_sub[24] ),
    .S(_02133_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__mux2_2 _29510_ (.A0(_02159_),
    .A1(\alu_add_sub[25] ),
    .S(_02133_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__mux2_2 _29511_ (.A0(_02160_),
    .A1(\alu_add_sub[26] ),
    .S(_02133_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__mux2_1 _29512_ (.A0(_02161_),
    .A1(\alu_add_sub[27] ),
    .S(_02133_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__mux2_2 _29513_ (.A0(_02162_),
    .A1(\alu_add_sub[28] ),
    .S(_02133_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__mux2_2 _29514_ (.A0(_02163_),
    .A1(\alu_add_sub[29] ),
    .S(_02133_),
    .X(\alu_out[29] ));
 sky130_fd_sc_hd__mux2_2 _29515_ (.A0(_02164_),
    .A1(\alu_add_sub[30] ),
    .S(_02133_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__mux2_2 _29516_ (.A0(_02165_),
    .A1(\alu_add_sub[31] ),
    .S(_02133_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__mux2_2 _29517_ (.A0(_02071_),
    .A1(\reg_next_pc[0] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[0] ));
 sky130_fd_sc_hd__mux2_4 _29518_ (.A0(_02072_),
    .A1(\reg_pc[1] ),
    .S(net439),
    .X(\cpuregs_wrdata[1] ));
 sky130_fd_sc_hd__mux2_2 _29519_ (.A0(_02074_),
    .A1(_02073_),
    .S(net439),
    .X(\cpuregs_wrdata[2] ));
 sky130_fd_sc_hd__mux2_2 _29520_ (.A0(_02076_),
    .A1(_02075_),
    .S(net439),
    .X(\cpuregs_wrdata[3] ));
 sky130_fd_sc_hd__mux2_2 _29521_ (.A0(_02078_),
    .A1(_02077_),
    .S(net439),
    .X(\cpuregs_wrdata[4] ));
 sky130_fd_sc_hd__mux2_2 _29522_ (.A0(_02080_),
    .A1(_02079_),
    .S(net439),
    .X(\cpuregs_wrdata[5] ));
 sky130_fd_sc_hd__mux2_2 _29523_ (.A0(_02082_),
    .A1(_02081_),
    .S(net439),
    .X(\cpuregs_wrdata[6] ));
 sky130_fd_sc_hd__mux2_4 _29524_ (.A0(_02084_),
    .A1(_02083_),
    .S(net439),
    .X(\cpuregs_wrdata[7] ));
 sky130_fd_sc_hd__mux2_4 _29525_ (.A0(_02086_),
    .A1(_02085_),
    .S(net439),
    .X(\cpuregs_wrdata[8] ));
 sky130_fd_sc_hd__mux2_4 _29526_ (.A0(_02088_),
    .A1(_02087_),
    .S(net439),
    .X(\cpuregs_wrdata[9] ));
 sky130_fd_sc_hd__mux2_4 _29527_ (.A0(_02090_),
    .A1(_02089_),
    .S(net439),
    .X(\cpuregs_wrdata[10] ));
 sky130_fd_sc_hd__mux2_4 _29528_ (.A0(_02092_),
    .A1(_02091_),
    .S(net439),
    .X(\cpuregs_wrdata[11] ));
 sky130_fd_sc_hd__mux2_4 _29529_ (.A0(_02094_),
    .A1(_02093_),
    .S(net439),
    .X(\cpuregs_wrdata[12] ));
 sky130_fd_sc_hd__mux2_2 _29530_ (.A0(_02096_),
    .A1(_02095_),
    .S(net439),
    .X(\cpuregs_wrdata[13] ));
 sky130_fd_sc_hd__mux2_4 _29531_ (.A0(_02098_),
    .A1(_02097_),
    .S(net439),
    .X(\cpuregs_wrdata[14] ));
 sky130_fd_sc_hd__mux2_4 _29532_ (.A0(_02100_),
    .A1(_02099_),
    .S(net439),
    .X(\cpuregs_wrdata[15] ));
 sky130_fd_sc_hd__mux2_4 _29533_ (.A0(_02102_),
    .A1(_02101_),
    .S(net439),
    .X(\cpuregs_wrdata[16] ));
 sky130_fd_sc_hd__mux2_2 _29534_ (.A0(_02104_),
    .A1(_02103_),
    .S(net439),
    .X(\cpuregs_wrdata[17] ));
 sky130_fd_sc_hd__mux2_4 _29535_ (.A0(_02106_),
    .A1(_02105_),
    .S(net439),
    .X(\cpuregs_wrdata[18] ));
 sky130_fd_sc_hd__mux2_4 _29536_ (.A0(_02108_),
    .A1(_02107_),
    .S(net439),
    .X(\cpuregs_wrdata[19] ));
 sky130_fd_sc_hd__mux2_2 _29537_ (.A0(_02110_),
    .A1(_02109_),
    .S(net439),
    .X(\cpuregs_wrdata[20] ));
 sky130_fd_sc_hd__mux2_4 _29538_ (.A0(_02112_),
    .A1(_02111_),
    .S(net439),
    .X(\cpuregs_wrdata[21] ));
 sky130_fd_sc_hd__mux2_4 _29539_ (.A0(_02114_),
    .A1(_02113_),
    .S(net439),
    .X(\cpuregs_wrdata[22] ));
 sky130_fd_sc_hd__mux2_4 _29540_ (.A0(_02116_),
    .A1(_02115_),
    .S(net439),
    .X(\cpuregs_wrdata[23] ));
 sky130_fd_sc_hd__mux2_4 _29541_ (.A0(_02118_),
    .A1(_02117_),
    .S(net439),
    .X(\cpuregs_wrdata[24] ));
 sky130_fd_sc_hd__mux2_2 _29542_ (.A0(_02120_),
    .A1(_02119_),
    .S(net439),
    .X(\cpuregs_wrdata[25] ));
 sky130_fd_sc_hd__mux2_4 _29543_ (.A0(_02122_),
    .A1(_02121_),
    .S(net439),
    .X(\cpuregs_wrdata[26] ));
 sky130_fd_sc_hd__mux2_4 _29544_ (.A0(_02124_),
    .A1(_02123_),
    .S(net439),
    .X(\cpuregs_wrdata[27] ));
 sky130_fd_sc_hd__mux2_4 _29545_ (.A0(_02126_),
    .A1(_02125_),
    .S(net439),
    .X(\cpuregs_wrdata[28] ));
 sky130_fd_sc_hd__mux2_4 _29546_ (.A0(_02128_),
    .A1(_02127_),
    .S(net439),
    .X(\cpuregs_wrdata[29] ));
 sky130_fd_sc_hd__mux2_4 _29547_ (.A0(_02130_),
    .A1(_02129_),
    .S(_02069_),
    .X(\cpuregs_wrdata[30] ));
 sky130_fd_sc_hd__mux2_4 _29548_ (.A0(_02132_),
    .A1(_02131_),
    .S(net439),
    .X(\cpuregs_wrdata[31] ));
 sky130_fd_sc_hd__mux2_1 _29549_ (.A0(_02316_),
    .A1(_02317_),
    .S(_00307_),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _29550_ (.A0(_00347_),
    .A1(_15210_),
    .S(_00336_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _29551_ (.A0(_15210_),
    .A1(_00348_),
    .S(net101),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _29552_ (.A0(_02304_),
    .A1(_02305_),
    .S(\irq_state[1] ),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _29553_ (.A0(_02306_),
    .A1(_02304_),
    .S(_02217_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _29554_ (.A0(_02214_),
    .A1(_02215_),
    .S(\irq_state[1] ),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _29555_ (.A0(_02216_),
    .A1(_02214_),
    .S(_02217_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _29556_ (.A0(_02218_),
    .A1(_02219_),
    .S(\irq_state[1] ),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _29557_ (.A0(_02220_),
    .A1(_02218_),
    .S(_02217_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _29558_ (.A0(_02221_),
    .A1(_02222_),
    .S(\irq_state[1] ),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _29559_ (.A0(_02223_),
    .A1(_02221_),
    .S(net421),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _29560_ (.A0(_02224_),
    .A1(_02225_),
    .S(\irq_state[1] ),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _29561_ (.A0(_02226_),
    .A1(_02224_),
    .S(net421),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _29562_ (.A0(_02227_),
    .A1(_02228_),
    .S(\irq_state[1] ),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _29563_ (.A0(_02229_),
    .A1(_02227_),
    .S(_02217_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _29564_ (.A0(_02230_),
    .A1(_02231_),
    .S(\irq_state[1] ),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _29565_ (.A0(_02232_),
    .A1(_02230_),
    .S(net421),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _29566_ (.A0(_02233_),
    .A1(_02234_),
    .S(\irq_state[1] ),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _29567_ (.A0(_02235_),
    .A1(_02233_),
    .S(net421),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _29568_ (.A0(_02236_),
    .A1(_02237_),
    .S(\irq_state[1] ),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _29569_ (.A0(_02238_),
    .A1(_02236_),
    .S(_02217_),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _29570_ (.A0(_02239_),
    .A1(_02240_),
    .S(\irq_state[1] ),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _29571_ (.A0(_02241_),
    .A1(_02239_),
    .S(net421),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _29572_ (.A0(_02242_),
    .A1(_02243_),
    .S(\irq_state[1] ),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _29573_ (.A0(_02244_),
    .A1(_02242_),
    .S(net421),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _29574_ (.A0(_02245_),
    .A1(_02246_),
    .S(\irq_state[1] ),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _29575_ (.A0(_02247_),
    .A1(_02245_),
    .S(net421),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _29576_ (.A0(_02248_),
    .A1(_02249_),
    .S(\irq_state[1] ),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _29577_ (.A0(_02250_),
    .A1(_02248_),
    .S(net421),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _29578_ (.A0(_02251_),
    .A1(_02252_),
    .S(\irq_state[1] ),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _29579_ (.A0(_02253_),
    .A1(_02251_),
    .S(net421),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _29580_ (.A0(_02254_),
    .A1(_02255_),
    .S(\irq_state[1] ),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _29581_ (.A0(_02256_),
    .A1(_02254_),
    .S(net421),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _29582_ (.A0(_02257_),
    .A1(_02258_),
    .S(\irq_state[1] ),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _29583_ (.A0(_02259_),
    .A1(_02257_),
    .S(net421),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _29584_ (.A0(_02260_),
    .A1(_02261_),
    .S(\irq_state[1] ),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _29585_ (.A0(_02262_),
    .A1(_02260_),
    .S(net421),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _29586_ (.A0(_02263_),
    .A1(_02264_),
    .S(\irq_state[1] ),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _29587_ (.A0(_02265_),
    .A1(_02263_),
    .S(net421),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _29588_ (.A0(_02266_),
    .A1(_02267_),
    .S(\irq_state[1] ),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _29589_ (.A0(_02268_),
    .A1(_02266_),
    .S(net421),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _29590_ (.A0(_02269_),
    .A1(_02270_),
    .S(\irq_state[1] ),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _29591_ (.A0(_02271_),
    .A1(_02269_),
    .S(net421),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _29592_ (.A0(_02272_),
    .A1(_02273_),
    .S(\irq_state[1] ),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _29593_ (.A0(_02274_),
    .A1(_02272_),
    .S(net421),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _29594_ (.A0(_02275_),
    .A1(_02276_),
    .S(\irq_state[1] ),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _29595_ (.A0(_02277_),
    .A1(_02275_),
    .S(net421),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _29596_ (.A0(_02278_),
    .A1(_02279_),
    .S(\irq_state[1] ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _29597_ (.A0(_02280_),
    .A1(_02278_),
    .S(net421),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _29598_ (.A0(_02281_),
    .A1(_02282_),
    .S(\irq_state[1] ),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _29599_ (.A0(_02283_),
    .A1(_02281_),
    .S(net421),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _29600_ (.A0(_02284_),
    .A1(_02285_),
    .S(\irq_state[1] ),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _29601_ (.A0(_02286_),
    .A1(_02284_),
    .S(net421),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _29602_ (.A0(_02287_),
    .A1(_02288_),
    .S(\irq_state[1] ),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _29603_ (.A0(_02289_),
    .A1(_02287_),
    .S(net421),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _29604_ (.A0(_02290_),
    .A1(_02291_),
    .S(\irq_state[1] ),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _29605_ (.A0(_02292_),
    .A1(_02290_),
    .S(net421),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _29606_ (.A0(_02293_),
    .A1(_02294_),
    .S(\irq_state[1] ),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _29607_ (.A0(_02295_),
    .A1(_02293_),
    .S(net421),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _29608_ (.A0(_02296_),
    .A1(_02297_),
    .S(\irq_state[1] ),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _29609_ (.A0(_02298_),
    .A1(_02296_),
    .S(net421),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _29610_ (.A0(_02299_),
    .A1(_02300_),
    .S(\irq_state[1] ),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _29611_ (.A0(_02301_),
    .A1(_02299_),
    .S(_02217_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_4 _29612_ (.A0(_01467_),
    .A1(\reg_next_pc[1] ),
    .S(_00292_),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_2 _29613_ (.A0(_00295_),
    .A1(\reg_next_pc[2] ),
    .S(_00292_),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_2 _29614_ (.A0(_01470_),
    .A1(\reg_next_pc[3] ),
    .S(net455),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_2 _29615_ (.A0(_01478_),
    .A1(\reg_next_pc[5] ),
    .S(net455),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_2 _29616_ (.A0(_01481_),
    .A1(\reg_next_pc[6] ),
    .S(net455),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_2 _29617_ (.A0(_01484_),
    .A1(\reg_next_pc[7] ),
    .S(net455),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_2 _29618_ (.A0(_01487_),
    .A1(\reg_next_pc[8] ),
    .S(net455),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_2 _29619_ (.A0(_01490_),
    .A1(\reg_next_pc[9] ),
    .S(net455),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_2 _29620_ (.A0(_01493_),
    .A1(\reg_next_pc[10] ),
    .S(net455),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_2 _29621_ (.A0(_01496_),
    .A1(\reg_next_pc[11] ),
    .S(net455),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_2 _29622_ (.A0(_01499_),
    .A1(\reg_next_pc[12] ),
    .S(net455),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_2 _29623_ (.A0(_01502_),
    .A1(\reg_next_pc[13] ),
    .S(net455),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_4 _29624_ (.A0(_01505_),
    .A1(\reg_next_pc[14] ),
    .S(net455),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_2 _29625_ (.A0(_01508_),
    .A1(\reg_next_pc[15] ),
    .S(net455),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_4 _29626_ (.A0(_01511_),
    .A1(\reg_next_pc[16] ),
    .S(net455),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_2 _29627_ (.A0(_01514_),
    .A1(\reg_next_pc[17] ),
    .S(net454),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_2 _29628_ (.A0(_01517_),
    .A1(\reg_next_pc[18] ),
    .S(net454),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_4 _29629_ (.A0(_01520_),
    .A1(\reg_next_pc[19] ),
    .S(net454),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_4 _29630_ (.A0(_01523_),
    .A1(\reg_next_pc[20] ),
    .S(net454),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_4 _29631_ (.A0(_01526_),
    .A1(\reg_next_pc[21] ),
    .S(net454),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_4 _29632_ (.A0(_01529_),
    .A1(\reg_next_pc[22] ),
    .S(net454),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_4 _29633_ (.A0(_01532_),
    .A1(\reg_next_pc[23] ),
    .S(net454),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_4 _29634_ (.A0(_01535_),
    .A1(\reg_next_pc[24] ),
    .S(net454),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_4 _29635_ (.A0(_01538_),
    .A1(\reg_next_pc[25] ),
    .S(net454),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_4 _29636_ (.A0(_01541_),
    .A1(\reg_next_pc[26] ),
    .S(net454),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_4 _29637_ (.A0(_01544_),
    .A1(\reg_next_pc[27] ),
    .S(net454),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_4 _29638_ (.A0(_01547_),
    .A1(\reg_next_pc[28] ),
    .S(net454),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_4 _29639_ (.A0(_01550_),
    .A1(\reg_next_pc[29] ),
    .S(net454),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_4 _29640_ (.A0(_01553_),
    .A1(\reg_next_pc[30] ),
    .S(net454),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_4 _29641_ (.A0(_01556_),
    .A1(\reg_next_pc[31] ),
    .S(_00292_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _29642_ (.A0(_00057_),
    .A1(_00064_),
    .S(net489),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _29643_ (.A0(_00065_),
    .A1(_02543_),
    .S(net488),
    .X(_15246_));
 sky130_fd_sc_hd__mux2_1 _29644_ (.A0(_00075_),
    .A1(_00082_),
    .S(net489),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _29645_ (.A0(_00083_),
    .A1(_02544_),
    .S(net488),
    .X(_15247_));
 sky130_fd_sc_hd__mux2_1 _29646_ (.A0(_00089_),
    .A1(_00092_),
    .S(net489),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _29647_ (.A0(_00093_),
    .A1(_02545_),
    .S(net488),
    .X(_15248_));
 sky130_fd_sc_hd__mux2_1 _29648_ (.A0(_00099_),
    .A1(_00102_),
    .S(net489),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _29649_ (.A0(_00103_),
    .A1(_02546_),
    .S(net488),
    .X(_15249_));
 sky130_fd_sc_hd__mux2_1 _29650_ (.A0(_00107_),
    .A1(_00108_),
    .S(net489),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _29651_ (.A0(_00109_),
    .A1(_02547_),
    .S(net488),
    .X(_15250_));
 sky130_fd_sc_hd__mux2_1 _29652_ (.A0(_00113_),
    .A1(_00114_),
    .S(net489),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _29653_ (.A0(_00115_),
    .A1(_02548_),
    .S(net488),
    .X(_15251_));
 sky130_fd_sc_hd__mux2_1 _29654_ (.A0(_00119_),
    .A1(_00120_),
    .S(net489),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _29655_ (.A0(_00121_),
    .A1(_02549_),
    .S(net488),
    .X(_15252_));
 sky130_fd_sc_hd__mux2_1 _29656_ (.A0(_00125_),
    .A1(_00126_),
    .S(net489),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _29657_ (.A0(_00127_),
    .A1(_02550_),
    .S(net488),
    .X(_15253_));
 sky130_fd_sc_hd__mux2_1 _29658_ (.A0(_00129_),
    .A1(_00106_),
    .S(net490),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _29659_ (.A0(_00130_),
    .A1(_00057_),
    .S(net489),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _29660_ (.A0(_00131_),
    .A1(_02551_),
    .S(net488),
    .X(_15254_));
 sky130_fd_sc_hd__mux2_1 _29661_ (.A0(_00133_),
    .A1(_00112_),
    .S(net490),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _29662_ (.A0(_00134_),
    .A1(_00075_),
    .S(net489),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _29663_ (.A0(_00135_),
    .A1(_02552_),
    .S(net488),
    .X(_15255_));
 sky130_fd_sc_hd__mux2_1 _29664_ (.A0(_00137_),
    .A1(_00118_),
    .S(net490),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _29665_ (.A0(_00138_),
    .A1(_00089_),
    .S(net489),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _29666_ (.A0(_00139_),
    .A1(_02553_),
    .S(net488),
    .X(_15256_));
 sky130_fd_sc_hd__mux2_1 _29667_ (.A0(_00141_),
    .A1(_00124_),
    .S(net490),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _29668_ (.A0(_00142_),
    .A1(_00099_),
    .S(net489),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _29669_ (.A0(_00143_),
    .A1(_02554_),
    .S(net488),
    .X(_15257_));
 sky130_fd_sc_hd__mux2_1 _29670_ (.A0(_00144_),
    .A1(_00136_),
    .S(net491),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _29671_ (.A0(_00145_),
    .A1(_00129_),
    .S(net490),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _29672_ (.A0(_00146_),
    .A1(_00107_),
    .S(net489),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _29673_ (.A0(_00147_),
    .A1(_02555_),
    .S(net488),
    .X(_15258_));
 sky130_fd_sc_hd__mux2_1 _29674_ (.A0(_00148_),
    .A1(_00140_),
    .S(net491),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _29675_ (.A0(_00149_),
    .A1(_00133_),
    .S(net490),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _29676_ (.A0(_00150_),
    .A1(_00113_),
    .S(net489),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _29677_ (.A0(_00151_),
    .A1(_02556_),
    .S(net488),
    .X(_15259_));
 sky130_fd_sc_hd__mux2_1 _29678_ (.A0(net329),
    .A1(net327),
    .S(net493),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _29679_ (.A0(_00152_),
    .A1(_00144_),
    .S(net491),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _29680_ (.A0(_00153_),
    .A1(_00137_),
    .S(net490),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _29681_ (.A0(_00154_),
    .A1(_00119_),
    .S(net489),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_2 _29682_ (.A0(_00155_),
    .A1(_02557_),
    .S(net488),
    .X(_15260_));
 sky130_fd_sc_hd__mux2_1 _29683_ (.A0(net330),
    .A1(net329),
    .S(net493),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _29684_ (.A0(_00156_),
    .A1(_00148_),
    .S(net491),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _29685_ (.A0(_00157_),
    .A1(_00141_),
    .S(net490),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _29686_ (.A0(_00158_),
    .A1(_00125_),
    .S(net489),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _29687_ (.A0(_00159_),
    .A1(_02558_),
    .S(net488),
    .X(_15261_));
 sky130_fd_sc_hd__mux2_1 _29688_ (.A0(net306),
    .A1(net317),
    .S(net200),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _29689_ (.A0(_00160_),
    .A1(_00161_),
    .S(net492),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _29690_ (.A0(_00162_),
    .A1(_00165_),
    .S(net490),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _29691_ (.A0(_00166_),
    .A1(_00173_),
    .S(net489),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _29692_ (.A0(_00174_),
    .A1(_00189_),
    .S(net488),
    .X(_15262_));
 sky130_fd_sc_hd__mux2_1 _29693_ (.A0(net317),
    .A1(net328),
    .S(net200),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _29694_ (.A0(_00190_),
    .A1(_00191_),
    .S(net492),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _29695_ (.A0(_00192_),
    .A1(_00195_),
    .S(net222),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _29696_ (.A0(_00196_),
    .A1(_00203_),
    .S(net225),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _29697_ (.A0(_00204_),
    .A1(_00220_),
    .S(net488),
    .X(_15273_));
 sky130_fd_sc_hd__mux2_1 _29698_ (.A0(_00161_),
    .A1(_00163_),
    .S(net492),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _29699_ (.A0(_00221_),
    .A1(_00222_),
    .S(net490),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _29700_ (.A0(_00223_),
    .A1(_00226_),
    .S(net489),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _29701_ (.A0(_00227_),
    .A1(_00234_),
    .S(net488),
    .X(_15284_));
 sky130_fd_sc_hd__mux2_1 _29702_ (.A0(_00191_),
    .A1(_00193_),
    .S(net492),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _29703_ (.A0(_00235_),
    .A1(_00236_),
    .S(net222),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _29704_ (.A0(_00237_),
    .A1(_00240_),
    .S(net489),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _29705_ (.A0(_00241_),
    .A1(_00248_),
    .S(net488),
    .X(_15287_));
 sky130_fd_sc_hd__mux2_1 _29706_ (.A0(_00165_),
    .A1(_00169_),
    .S(net490),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _29707_ (.A0(_00249_),
    .A1(_00250_),
    .S(net489),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _29708_ (.A0(_00251_),
    .A1(_00254_),
    .S(net488),
    .X(_15288_));
 sky130_fd_sc_hd__mux2_1 _29709_ (.A0(_00195_),
    .A1(_00199_),
    .S(net222),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _29710_ (.A0(_00255_),
    .A1(_00256_),
    .S(net225),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _29711_ (.A0(_00257_),
    .A1(_00260_),
    .S(net488),
    .X(_15289_));
 sky130_fd_sc_hd__mux2_1 _29712_ (.A0(_00222_),
    .A1(_00224_),
    .S(net490),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _29713_ (.A0(_00261_),
    .A1(_00262_),
    .S(net489),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _29714_ (.A0(_00263_),
    .A1(_00266_),
    .S(net488),
    .X(_15290_));
 sky130_fd_sc_hd__mux2_1 _29715_ (.A0(_00236_),
    .A1(_00238_),
    .S(net222),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _29716_ (.A0(_00267_),
    .A1(_00268_),
    .S(net225),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _29717_ (.A0(_00269_),
    .A1(_00272_),
    .S(net488),
    .X(_15291_));
 sky130_fd_sc_hd__mux2_1 _29718_ (.A0(_00173_),
    .A1(_00181_),
    .S(net489),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _29719_ (.A0(_00273_),
    .A1(_00274_),
    .S(net488),
    .X(_15292_));
 sky130_fd_sc_hd__mux2_1 _29720_ (.A0(_00203_),
    .A1(_00211_),
    .S(net225),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _29721_ (.A0(_00275_),
    .A1(_00276_),
    .S(net488),
    .X(_15293_));
 sky130_fd_sc_hd__mux2_1 _29722_ (.A0(_00226_),
    .A1(_00230_),
    .S(net489),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _29723_ (.A0(_00277_),
    .A1(_00278_),
    .S(net488),
    .X(_15263_));
 sky130_fd_sc_hd__mux2_1 _29724_ (.A0(_00240_),
    .A1(_00244_),
    .S(net225),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _29725_ (.A0(_00279_),
    .A1(_00280_),
    .S(net488),
    .X(_15264_));
 sky130_fd_sc_hd__mux2_1 _29726_ (.A0(_00250_),
    .A1(_00252_),
    .S(net489),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _29727_ (.A0(_00281_),
    .A1(_00282_),
    .S(net488),
    .X(_15265_));
 sky130_fd_sc_hd__mux2_1 _29728_ (.A0(_00256_),
    .A1(_00258_),
    .S(net225),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _29729_ (.A0(_00283_),
    .A1(_00284_),
    .S(net226),
    .X(_15266_));
 sky130_fd_sc_hd__mux2_1 _29730_ (.A0(_00262_),
    .A1(_00264_),
    .S(net489),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _29731_ (.A0(_00285_),
    .A1(_00286_),
    .S(net488),
    .X(_15267_));
 sky130_fd_sc_hd__mux2_1 _29732_ (.A0(_00268_),
    .A1(_00270_),
    .S(net225),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _29733_ (.A0(_00287_),
    .A1(_00288_),
    .S(net226),
    .X(_15268_));
 sky130_fd_sc_hd__mux2_1 _29734_ (.A0(_00189_),
    .A1(_00216_),
    .S(net488),
    .X(_15269_));
 sky130_fd_sc_hd__mux2_1 _29735_ (.A0(_00220_),
    .A1(_00216_),
    .S(net488),
    .X(_15270_));
 sky130_fd_sc_hd__mux2_1 _29736_ (.A0(_00234_),
    .A1(_00216_),
    .S(net488),
    .X(_15271_));
 sky130_fd_sc_hd__mux2_1 _29737_ (.A0(_00248_),
    .A1(_00216_),
    .S(net226),
    .X(_15272_));
 sky130_fd_sc_hd__mux2_1 _29738_ (.A0(_00254_),
    .A1(_00216_),
    .S(net488),
    .X(_15274_));
 sky130_fd_sc_hd__mux2_1 _29739_ (.A0(_00260_),
    .A1(_00216_),
    .S(net226),
    .X(_15275_));
 sky130_fd_sc_hd__mux2_1 _29740_ (.A0(_00266_),
    .A1(_00216_),
    .S(net488),
    .X(_15276_));
 sky130_fd_sc_hd__mux2_1 _29741_ (.A0(_00272_),
    .A1(_00216_),
    .S(net226),
    .X(_15277_));
 sky130_fd_sc_hd__mux2_1 _29742_ (.A0(_00274_),
    .A1(_00216_),
    .S(net488),
    .X(_15278_));
 sky130_fd_sc_hd__mux2_1 _29743_ (.A0(_00276_),
    .A1(_00216_),
    .S(net488),
    .X(_15279_));
 sky130_fd_sc_hd__mux2_1 _29744_ (.A0(_00278_),
    .A1(_00216_),
    .S(net488),
    .X(_15280_));
 sky130_fd_sc_hd__mux2_1 _29745_ (.A0(_00280_),
    .A1(_00216_),
    .S(net488),
    .X(_15281_));
 sky130_fd_sc_hd__mux2_1 _29746_ (.A0(_00282_),
    .A1(_00216_),
    .S(net488),
    .X(_15282_));
 sky130_fd_sc_hd__mux2_1 _29747_ (.A0(_00284_),
    .A1(_00216_),
    .S(net226),
    .X(_15283_));
 sky130_fd_sc_hd__mux2_1 _29748_ (.A0(_00286_),
    .A1(_00216_),
    .S(net488),
    .X(_15285_));
 sky130_fd_sc_hd__mux2_1 _29749_ (.A0(_00288_),
    .A1(_00216_),
    .S(net226),
    .X(_15286_));
 sky130_fd_sc_hd__mux2_1 _29750_ (.A0(_01697_),
    .A1(_01698_),
    .S(\irq_state[1] ),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _29751_ (.A0(_01705_),
    .A1(_01699_),
    .S(_01700_),
    .X(_15245_));
 sky130_fd_sc_hd__mux2_1 _29752_ (.A0(_01720_),
    .A1(\irq_pending[0] ),
    .S(_01706_),
    .X(_15211_));
 sky130_fd_sc_hd__mux2_1 _29753_ (.A0(_01733_),
    .A1(\irq_pending[1] ),
    .S(_01706_),
    .X(_15222_));
 sky130_fd_sc_hd__mux2_1 _29754_ (.A0(_01746_),
    .A1(\irq_pending[2] ),
    .S(_01706_),
    .X(_15233_));
 sky130_fd_sc_hd__mux2_1 _29755_ (.A0(_01759_),
    .A1(\irq_pending[3] ),
    .S(_01706_),
    .X(_15236_));
 sky130_fd_sc_hd__mux2_1 _29756_ (.A0(_01772_),
    .A1(\irq_pending[4] ),
    .S(_01706_),
    .X(_15237_));
 sky130_fd_sc_hd__mux2_1 _29757_ (.A0(_01785_),
    .A1(\irq_pending[5] ),
    .S(_01706_),
    .X(_15238_));
 sky130_fd_sc_hd__mux2_1 _29758_ (.A0(_01798_),
    .A1(\irq_pending[6] ),
    .S(_01706_),
    .X(_15239_));
 sky130_fd_sc_hd__mux2_1 _29759_ (.A0(_01811_),
    .A1(\irq_pending[7] ),
    .S(_01706_),
    .X(_15240_));
 sky130_fd_sc_hd__mux2_2 _29760_ (.A0(_01825_),
    .A1(\irq_pending[8] ),
    .S(_01706_),
    .X(_15241_));
 sky130_fd_sc_hd__mux2_1 _29761_ (.A0(_01838_),
    .A1(\irq_pending[9] ),
    .S(net436),
    .X(_15242_));
 sky130_fd_sc_hd__mux2_2 _29762_ (.A0(_01851_),
    .A1(\irq_pending[10] ),
    .S(_01706_),
    .X(_15212_));
 sky130_fd_sc_hd__mux2_2 _29763_ (.A0(_01864_),
    .A1(\irq_pending[11] ),
    .S(net436),
    .X(_15213_));
 sky130_fd_sc_hd__mux2_2 _29764_ (.A0(_01877_),
    .A1(\irq_pending[12] ),
    .S(_01706_),
    .X(_15214_));
 sky130_fd_sc_hd__mux2_1 _29765_ (.A0(_01890_),
    .A1(\irq_pending[13] ),
    .S(net436),
    .X(_15215_));
 sky130_fd_sc_hd__mux2_1 _29766_ (.A0(_01903_),
    .A1(\irq_pending[14] ),
    .S(net436),
    .X(_15216_));
 sky130_fd_sc_hd__mux2_2 _29767_ (.A0(_01916_),
    .A1(\irq_pending[15] ),
    .S(net436),
    .X(_15217_));
 sky130_fd_sc_hd__mux2_1 _29768_ (.A0(_01925_),
    .A1(\irq_pending[16] ),
    .S(net436),
    .X(_15218_));
 sky130_fd_sc_hd__mux2_1 _29769_ (.A0(_01934_),
    .A1(\irq_pending[17] ),
    .S(net436),
    .X(_15219_));
 sky130_fd_sc_hd__mux2_1 _29770_ (.A0(_01943_),
    .A1(\irq_pending[18] ),
    .S(net436),
    .X(_15220_));
 sky130_fd_sc_hd__mux2_1 _29771_ (.A0(_01952_),
    .A1(\irq_pending[19] ),
    .S(net436),
    .X(_15221_));
 sky130_fd_sc_hd__mux2_1 _29772_ (.A0(_01961_),
    .A1(\irq_pending[20] ),
    .S(net436),
    .X(_15223_));
 sky130_fd_sc_hd__mux2_1 _29773_ (.A0(_01970_),
    .A1(\irq_pending[21] ),
    .S(net436),
    .X(_15224_));
 sky130_fd_sc_hd__mux2_1 _29774_ (.A0(_01979_),
    .A1(\irq_pending[22] ),
    .S(net436),
    .X(_15225_));
 sky130_fd_sc_hd__mux2_1 _29775_ (.A0(_01988_),
    .A1(\irq_pending[23] ),
    .S(net436),
    .X(_15226_));
 sky130_fd_sc_hd__mux2_1 _29776_ (.A0(_01997_),
    .A1(\irq_pending[24] ),
    .S(net436),
    .X(_15227_));
 sky130_fd_sc_hd__mux2_1 _29777_ (.A0(_02006_),
    .A1(\irq_pending[25] ),
    .S(net436),
    .X(_15228_));
 sky130_fd_sc_hd__mux2_1 _29778_ (.A0(_02015_),
    .A1(\irq_pending[26] ),
    .S(net436),
    .X(_15229_));
 sky130_fd_sc_hd__mux2_1 _29779_ (.A0(_02024_),
    .A1(\irq_pending[27] ),
    .S(_01706_),
    .X(_15230_));
 sky130_fd_sc_hd__mux2_1 _29780_ (.A0(_02033_),
    .A1(\irq_pending[28] ),
    .S(net436),
    .X(_15231_));
 sky130_fd_sc_hd__mux2_1 _29781_ (.A0(_02042_),
    .A1(\irq_pending[29] ),
    .S(_01706_),
    .X(_15232_));
 sky130_fd_sc_hd__mux2_1 _29782_ (.A0(_02051_),
    .A1(\irq_pending[30] ),
    .S(_01706_),
    .X(_15234_));
 sky130_fd_sc_hd__mux2_1 _29783_ (.A0(_02060_),
    .A1(\irq_pending[31] ),
    .S(net436),
    .X(_15235_));
 sky130_fd_sc_hd__mux2_1 _29784_ (.A0(_02061_),
    .A1(\cpu_state[2] ),
    .S(_02542_),
    .X(_15206_));
 sky130_fd_sc_hd__mux2_1 _29785_ (.A0(\decoded_rd[0] ),
    .A1(\irq_state[0] ),
    .S(_00308_),
    .X(_15205_));
 sky130_fd_sc_hd__mux2_1 _29786_ (.A0(_02062_),
    .A1(_02065_),
    .S(_02542_),
    .X(_15243_));
 sky130_fd_sc_hd__mux2_1 _29787_ (.A0(_02068_),
    .A1(_02066_),
    .S(_02067_),
    .X(_15244_));
 sky130_fd_sc_hd__mux2_1 _29788_ (.A0(_02166_),
    .A1(_00291_),
    .S(_00290_),
    .X(_15207_));
 sky130_fd_sc_hd__mux2_1 _29789_ (.A0(_02166_),
    .A1(mem_do_wdata),
    .S(_00290_),
    .X(_15208_));
 sky130_fd_sc_hd__mux2_1 _29790_ (.A0(_00271_),
    .A1(_00216_),
    .S(net225),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _29791_ (.A0(_00265_),
    .A1(_00216_),
    .S(net489),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _29792_ (.A0(_00259_),
    .A1(_00216_),
    .S(net225),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _29793_ (.A0(_00253_),
    .A1(_00216_),
    .S(net489),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _29794_ (.A0(_00247_),
    .A1(_00216_),
    .S(net225),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _29795_ (.A0(_00233_),
    .A1(_00216_),
    .S(net489),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _29796_ (.A0(_00219_),
    .A1(_00216_),
    .S(net225),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _29797_ (.A0(_00188_),
    .A1(_00216_),
    .S(net489),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _29798_ (.A0(_00270_),
    .A1(_00271_),
    .S(net225),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _29799_ (.A0(_00246_),
    .A1(_00216_),
    .S(net222),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _29800_ (.A0(_00243_),
    .A1(_00245_),
    .S(net222),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _29801_ (.A0(_00239_),
    .A1(_00242_),
    .S(net222),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _29802_ (.A0(_00264_),
    .A1(_00265_),
    .S(net489),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _29803_ (.A0(_00232_),
    .A1(_00216_),
    .S(net490),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _29804_ (.A0(_00229_),
    .A1(_00231_),
    .S(net490),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _29805_ (.A0(_00225_),
    .A1(_00228_),
    .S(net490),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _29806_ (.A0(_00258_),
    .A1(_00259_),
    .S(net225),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _29807_ (.A0(_00218_),
    .A1(_00216_),
    .S(net222),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _29808_ (.A0(_00210_),
    .A1(_00214_),
    .S(net222),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _29809_ (.A0(_00202_),
    .A1(_00207_),
    .S(net222),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _29810_ (.A0(_00252_),
    .A1(_00253_),
    .S(net489),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _29811_ (.A0(_00187_),
    .A1(_00216_),
    .S(net490),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _29812_ (.A0(_00180_),
    .A1(_00184_),
    .S(net490),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _29813_ (.A0(_00172_),
    .A1(_00177_),
    .S(net490),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _29814_ (.A0(_00244_),
    .A1(_00247_),
    .S(net225),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _29815_ (.A0(_00245_),
    .A1(_00246_),
    .S(net222),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _29816_ (.A0(_00217_),
    .A1(_00216_),
    .S(net492),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _29817_ (.A0(_00213_),
    .A1(_00215_),
    .S(net492),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _29818_ (.A0(_00242_),
    .A1(_00243_),
    .S(net222),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _29819_ (.A0(_00209_),
    .A1(_00212_),
    .S(net492),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _29820_ (.A0(_00206_),
    .A1(_00208_),
    .S(net492),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _29821_ (.A0(_00238_),
    .A1(_00239_),
    .S(net222),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _29822_ (.A0(_00201_),
    .A1(_00205_),
    .S(net492),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _29823_ (.A0(_00198_),
    .A1(_00200_),
    .S(net492),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _29824_ (.A0(_00194_),
    .A1(_00197_),
    .S(net492),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _29825_ (.A0(_00230_),
    .A1(_00233_),
    .S(net489),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _29826_ (.A0(_00231_),
    .A1(_00232_),
    .S(net490),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _29827_ (.A0(_00186_),
    .A1(_00216_),
    .S(net492),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _29828_ (.A0(_00183_),
    .A1(_00185_),
    .S(net492),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _29829_ (.A0(_00228_),
    .A1(_00229_),
    .S(net490),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _29830_ (.A0(_00179_),
    .A1(_00182_),
    .S(net492),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _29831_ (.A0(_00176_),
    .A1(_00178_),
    .S(net492),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _29832_ (.A0(_00224_),
    .A1(_00225_),
    .S(net490),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _29833_ (.A0(_00171_),
    .A1(_00175_),
    .S(net492),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _29834_ (.A0(_00168_),
    .A1(_00170_),
    .S(net492),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _29835_ (.A0(_00164_),
    .A1(_00167_),
    .S(net492),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _29836_ (.A0(_00211_),
    .A1(_00219_),
    .S(net225),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _29837_ (.A0(_00214_),
    .A1(_00218_),
    .S(net222),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _29838_ (.A0(_00215_),
    .A1(_00217_),
    .S(net492),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _29839_ (.A0(net330),
    .A1(_00216_),
    .S(net200),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _29840_ (.A0(net327),
    .A1(net329),
    .S(net200),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _29841_ (.A0(_00212_),
    .A1(_00213_),
    .S(net492),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _29842_ (.A0(net325),
    .A1(net326),
    .S(net200),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _29843_ (.A0(net323),
    .A1(net324),
    .S(net200),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _29844_ (.A0(_00207_),
    .A1(_00210_),
    .S(net222),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _29845_ (.A0(_00208_),
    .A1(_00209_),
    .S(net492),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _29846_ (.A0(net321),
    .A1(net322),
    .S(net200),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _29847_ (.A0(net319),
    .A1(net320),
    .S(net200),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _29848_ (.A0(_00205_),
    .A1(_00206_),
    .S(net492),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _29849_ (.A0(net316),
    .A1(net318),
    .S(net200),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _29850_ (.A0(net314),
    .A1(net315),
    .S(net200),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _29851_ (.A0(_00199_),
    .A1(_00202_),
    .S(net222),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _29852_ (.A0(_00200_),
    .A1(_00201_),
    .S(net492),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _29853_ (.A0(net312),
    .A1(net313),
    .S(net200),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _29854_ (.A0(net310),
    .A1(net311),
    .S(net200),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _29855_ (.A0(_00197_),
    .A1(_00198_),
    .S(net492),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _29856_ (.A0(net308),
    .A1(net309),
    .S(net200),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _29857_ (.A0(net337),
    .A1(net307),
    .S(net200),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _29858_ (.A0(_00193_),
    .A1(_00194_),
    .S(net492),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _29859_ (.A0(net335),
    .A1(net336),
    .S(net200),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _29860_ (.A0(net333),
    .A1(net334),
    .S(net200),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _29861_ (.A0(net331),
    .A1(net332),
    .S(net200),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _29862_ (.A0(_00181_),
    .A1(_00188_),
    .S(net489),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _29863_ (.A0(_00184_),
    .A1(_00187_),
    .S(net490),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _29864_ (.A0(_00185_),
    .A1(_00186_),
    .S(net492),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _29865_ (.A0(net329),
    .A1(net330),
    .S(net493),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _29866_ (.A0(net326),
    .A1(net327),
    .S(net493),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _29867_ (.A0(_00182_),
    .A1(_00183_),
    .S(net492),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _29868_ (.A0(net324),
    .A1(net325),
    .S(net493),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _29869_ (.A0(net322),
    .A1(net323),
    .S(net493),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _29870_ (.A0(_00177_),
    .A1(_00180_),
    .S(net490),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _29871_ (.A0(_00178_),
    .A1(_00179_),
    .S(net492),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _29872_ (.A0(net320),
    .A1(net321),
    .S(net493),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _29873_ (.A0(net318),
    .A1(net319),
    .S(net493),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _29874_ (.A0(_00175_),
    .A1(_00176_),
    .S(net492),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _29875_ (.A0(net315),
    .A1(net316),
    .S(net493),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _29876_ (.A0(net313),
    .A1(net314),
    .S(net493),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _29877_ (.A0(_00169_),
    .A1(_00172_),
    .S(net490),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _29878_ (.A0(_00170_),
    .A1(_00171_),
    .S(net492),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _29879_ (.A0(net311),
    .A1(net312),
    .S(net493),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _29880_ (.A0(net309),
    .A1(net310),
    .S(net493),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _29881_ (.A0(_00167_),
    .A1(_00168_),
    .S(net492),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _29882_ (.A0(net307),
    .A1(net308),
    .S(net493),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _29883_ (.A0(net336),
    .A1(net337),
    .S(net493),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _29884_ (.A0(_00163_),
    .A1(_00164_),
    .S(net492),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _29885_ (.A0(net334),
    .A1(net335),
    .S(net493),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _29886_ (.A0(net332),
    .A1(net333),
    .S(net493),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _29887_ (.A0(net328),
    .A1(net331),
    .S(net200),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _29888_ (.A0(net327),
    .A1(net326),
    .S(net493),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _29889_ (.A0(net326),
    .A1(net325),
    .S(net493),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _29890_ (.A0(_00140_),
    .A1(_00132_),
    .S(net491),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _29891_ (.A0(net325),
    .A1(net324),
    .S(net493),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _29892_ (.A0(_00136_),
    .A1(_00128_),
    .S(net491),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _29893_ (.A0(net324),
    .A1(net323),
    .S(net493),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _29894_ (.A0(_00132_),
    .A1(_00123_),
    .S(net491),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _29895_ (.A0(net323),
    .A1(net322),
    .S(net493),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _29896_ (.A0(_00128_),
    .A1(_00117_),
    .S(net491),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _29897_ (.A0(net322),
    .A1(net321),
    .S(net493),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _29898_ (.A0(_00098_),
    .A1(_00100_),
    .S(net490),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _29899_ (.A0(_00124_),
    .A1(_00097_),
    .S(net490),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _29900_ (.A0(_00123_),
    .A1(_00111_),
    .S(net491),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _29901_ (.A0(net321),
    .A1(net320),
    .S(net493),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _29902_ (.A0(_00101_),
    .A1(_00094_),
    .S(net490),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _29903_ (.A0(_00088_),
    .A1(_00090_),
    .S(net490),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _29904_ (.A0(_00118_),
    .A1(_00087_),
    .S(net490),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _29905_ (.A0(_00117_),
    .A1(_00105_),
    .S(net491),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _29906_ (.A0(net320),
    .A1(net319),
    .S(net493),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _29907_ (.A0(_00091_),
    .A1(_00084_),
    .S(net490),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _29908_ (.A0(_00074_),
    .A1(_00078_),
    .S(net490),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _29909_ (.A0(_00112_),
    .A1(_00071_),
    .S(net490),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _29910_ (.A0(_00111_),
    .A1(_00096_),
    .S(net491),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _29911_ (.A0(net319),
    .A1(net318),
    .S(net493),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _29912_ (.A0(_00081_),
    .A1(_00067_),
    .S(net490),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _29913_ (.A0(_00056_),
    .A1(_00060_),
    .S(net490),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _29914_ (.A0(_00106_),
    .A1(_00053_),
    .S(net490),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _29915_ (.A0(_00105_),
    .A1(_00086_),
    .S(net491),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _29916_ (.A0(net318),
    .A1(net316),
    .S(net493),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _29917_ (.A0(_00063_),
    .A1(_00049_),
    .S(net222),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _29918_ (.A0(_00100_),
    .A1(_00101_),
    .S(net490),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _29919_ (.A0(_00077_),
    .A1(_00079_),
    .S(net491),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _29920_ (.A0(_00073_),
    .A1(_00076_),
    .S(net491),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _29921_ (.A0(_00097_),
    .A1(_00098_),
    .S(net490),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _29922_ (.A0(_00070_),
    .A1(_00072_),
    .S(net491),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _29923_ (.A0(_00096_),
    .A1(_00069_),
    .S(net491),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _29924_ (.A0(net316),
    .A1(net315),
    .S(net493),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_2 _29925_ (.A0(_00080_),
    .A1(_00066_),
    .S(net491),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _29926_ (.A0(_00090_),
    .A1(_00091_),
    .S(net490),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _29927_ (.A0(_00059_),
    .A1(_00061_),
    .S(net491),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _29928_ (.A0(_00055_),
    .A1(_00058_),
    .S(net491),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _29929_ (.A0(_00087_),
    .A1(_00088_),
    .S(net490),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _29930_ (.A0(_00052_),
    .A1(_00054_),
    .S(net491),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _29931_ (.A0(_00086_),
    .A1(_00051_),
    .S(net491),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _29932_ (.A0(net315),
    .A1(net314),
    .S(net493),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_2 _29933_ (.A0(_00062_),
    .A1(_00048_),
    .S(net491),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _29934_ (.A0(_00078_),
    .A1(_00081_),
    .S(net490),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _29935_ (.A0(_00079_),
    .A1(_00080_),
    .S(net491),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _29936_ (.A0(net331),
    .A1(net328),
    .S(net200),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _29937_ (.A0(net333),
    .A1(net332),
    .S(net493),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _29938_ (.A0(_00076_),
    .A1(_00077_),
    .S(net491),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _29939_ (.A0(net335),
    .A1(net334),
    .S(net493),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _29940_ (.A0(net337),
    .A1(net336),
    .S(net493),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _29941_ (.A0(_00071_),
    .A1(_00074_),
    .S(net490),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _29942_ (.A0(_00072_),
    .A1(_00073_),
    .S(net491),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _29943_ (.A0(net308),
    .A1(net307),
    .S(net493),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _29944_ (.A0(net310),
    .A1(net309),
    .S(net493),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _29945_ (.A0(_00069_),
    .A1(_00070_),
    .S(net491),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _29946_ (.A0(net312),
    .A1(net311),
    .S(net493),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _29947_ (.A0(net314),
    .A1(net313),
    .S(net493),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_2 _29948_ (.A0(net317),
    .A1(net306),
    .S(net200),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _29949_ (.A0(_00060_),
    .A1(_00063_),
    .S(net490),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _29950_ (.A0(_00061_),
    .A1(_00062_),
    .S(net491),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _29951_ (.A0(net328),
    .A1(net317),
    .S(net200),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _29952_ (.A0(net332),
    .A1(net331),
    .S(net493),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _29953_ (.A0(_00058_),
    .A1(_00059_),
    .S(net491),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _29954_ (.A0(net334),
    .A1(net333),
    .S(net493),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _29955_ (.A0(net336),
    .A1(net335),
    .S(net493),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _29956_ (.A0(_00053_),
    .A1(_00056_),
    .S(net490),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _29957_ (.A0(_00054_),
    .A1(_00055_),
    .S(net491),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _29958_ (.A0(net307),
    .A1(net337),
    .S(net493),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _29959_ (.A0(net309),
    .A1(net308),
    .S(net493),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _29960_ (.A0(_00051_),
    .A1(_00052_),
    .S(net491),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _29961_ (.A0(net311),
    .A1(net310),
    .S(net493),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _29962_ (.A0(net313),
    .A1(net312),
    .S(net493),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _29963_ (.A0(_02408_),
    .A1(net362),
    .S(instr_sub),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_2 _29964_ (.A0(_02406_),
    .A1(_02405_),
    .S(instr_sub),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _29965_ (.A0(_02403_),
    .A1(_02402_),
    .S(instr_sub),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_2 _29966_ (.A0(_02400_),
    .A1(_02399_),
    .S(instr_sub),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_2 _29967_ (.A0(_02397_),
    .A1(_02396_),
    .S(instr_sub),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_2 _29968_ (.A0(_02394_),
    .A1(_02393_),
    .S(instr_sub),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_2 _29969_ (.A0(_02391_),
    .A1(_02390_),
    .S(instr_sub),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_2 _29970_ (.A0(_02388_),
    .A1(_02387_),
    .S(instr_sub),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _29971_ (.A0(_02385_),
    .A1(_02384_),
    .S(instr_sub),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _29972_ (.A0(_02382_),
    .A1(_02381_),
    .S(instr_sub),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _29973_ (.A0(_02379_),
    .A1(_02378_),
    .S(instr_sub),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_2 _29974_ (.A0(_02376_),
    .A1(_02375_),
    .S(instr_sub),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _29975_ (.A0(_02373_),
    .A1(_02372_),
    .S(instr_sub),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_2 _29976_ (.A0(_02370_),
    .A1(_02369_),
    .S(instr_sub),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_2 _29977_ (.A0(_02367_),
    .A1(_02366_),
    .S(instr_sub),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_2 _29978_ (.A0(_02364_),
    .A1(_02363_),
    .S(instr_sub),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_2 _29979_ (.A0(_02361_),
    .A1(_02360_),
    .S(instr_sub),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_2 _29980_ (.A0(_02358_),
    .A1(_02357_),
    .S(instr_sub),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_2 _29981_ (.A0(_02355_),
    .A1(_02354_),
    .S(instr_sub),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_2 _29982_ (.A0(_02352_),
    .A1(_02351_),
    .S(instr_sub),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_2 _29983_ (.A0(_02349_),
    .A1(_02348_),
    .S(instr_sub),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_2 _29984_ (.A0(_02346_),
    .A1(_02345_),
    .S(instr_sub),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_2 _29985_ (.A0(_02343_),
    .A1(_02342_),
    .S(instr_sub),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_2 _29986_ (.A0(_02340_),
    .A1(_02339_),
    .S(instr_sub),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_2 _29987_ (.A0(_02337_),
    .A1(_02336_),
    .S(instr_sub),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_2 _29988_ (.A0(_02334_),
    .A1(_02333_),
    .S(instr_sub),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _29989_ (.A0(_02331_),
    .A1(_02330_),
    .S(instr_sub),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _29990_ (.A0(_02328_),
    .A1(_02327_),
    .S(instr_sub),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _29991_ (.A0(_02325_),
    .A1(_02324_),
    .S(instr_sub),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _29992_ (.A0(_02322_),
    .A1(_02321_),
    .S(instr_sub),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_2 _29993_ (.A0(_02319_),
    .A1(_02318_),
    .S(instr_sub),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _29994_ (.A0(_02313_),
    .A1(_02314_),
    .S(_00306_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _29995_ (.A0(_02311_),
    .A1(_02315_),
    .S(_00303_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _29996_ (.A0(_02311_),
    .A1(_02312_),
    .S(_00305_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _29997_ (.A0(_02307_),
    .A1(_02308_),
    .S(\irq_state[1] ),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _29998_ (.A0(_02309_),
    .A1(_02307_),
    .S(_02217_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _29999_ (.A0(_02302_),
    .A1(\irq_pending[0] ),
    .S(net417),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _30000_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(latched_stalu),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _30001_ (.A0(_02063_),
    .A1(_00343_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _30002_ (.A0(_02056_),
    .A1(_02055_),
    .S(net485),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_2 _30003_ (.A0(_02058_),
    .A1(_02057_),
    .S(_01717_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _30004_ (.A0(\pcpi_mul.rd[31] ),
    .A1(\pcpi_mul.rd[63] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _30005_ (.A0(_01908_),
    .A1(_02052_),
    .S(_01816_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _30006_ (.A0(_02047_),
    .A1(_02046_),
    .S(net485),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _30007_ (.A0(_02049_),
    .A1(_02048_),
    .S(net446),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _30008_ (.A0(\pcpi_mul.rd[30] ),
    .A1(\pcpi_mul.rd[62] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _30009_ (.A0(_01908_),
    .A1(_02043_),
    .S(net481),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _30010_ (.A0(_02038_),
    .A1(_02037_),
    .S(net485),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_2 _30011_ (.A0(_02040_),
    .A1(_02039_),
    .S(_01717_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _30012_ (.A0(\pcpi_mul.rd[29] ),
    .A1(\pcpi_mul.rd[61] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _30013_ (.A0(_01908_),
    .A1(_02034_),
    .S(net481),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _30014_ (.A0(_02029_),
    .A1(_02028_),
    .S(_01714_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _30015_ (.A0(_02031_),
    .A1(_02030_),
    .S(_01717_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _30016_ (.A0(\pcpi_mul.rd[28] ),
    .A1(\pcpi_mul.rd[60] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _30017_ (.A0(_01908_),
    .A1(_02025_),
    .S(net481),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _30018_ (.A0(_02020_),
    .A1(_02019_),
    .S(net487),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_2 _30019_ (.A0(_02022_),
    .A1(_02021_),
    .S(net446),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _30020_ (.A0(\pcpi_mul.rd[27] ),
    .A1(\pcpi_mul.rd[59] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _30021_ (.A0(_01908_),
    .A1(_02016_),
    .S(net481),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _30022_ (.A0(_02011_),
    .A1(_02010_),
    .S(_01714_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_2 _30023_ (.A0(_02013_),
    .A1(_02012_),
    .S(_01717_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _30024_ (.A0(\pcpi_mul.rd[26] ),
    .A1(\pcpi_mul.rd[58] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _30025_ (.A0(_01908_),
    .A1(_02007_),
    .S(net481),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _30026_ (.A0(_02002_),
    .A1(_02001_),
    .S(_01714_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_2 _30027_ (.A0(_02004_),
    .A1(_02003_),
    .S(_01717_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_2 _30028_ (.A0(\pcpi_mul.rd[25] ),
    .A1(\pcpi_mul.rd[57] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _30029_ (.A0(_01908_),
    .A1(_01998_),
    .S(net481),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _30030_ (.A0(_01993_),
    .A1(_01992_),
    .S(net487),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _30031_ (.A0(_01995_),
    .A1(_01994_),
    .S(net446),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_2 _30032_ (.A0(\pcpi_mul.rd[24] ),
    .A1(\pcpi_mul.rd[56] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _30033_ (.A0(_01908_),
    .A1(_01989_),
    .S(net481),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _30034_ (.A0(_01984_),
    .A1(_01983_),
    .S(net487),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_2 _30035_ (.A0(_01986_),
    .A1(_01985_),
    .S(_01717_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_2 _30036_ (.A0(\pcpi_mul.rd[23] ),
    .A1(\pcpi_mul.rd[55] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _30037_ (.A0(_01908_),
    .A1(_01980_),
    .S(net481),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _30038_ (.A0(_01975_),
    .A1(_01974_),
    .S(_01714_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_2 _30039_ (.A0(_01977_),
    .A1(_01976_),
    .S(_01717_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_2 _30040_ (.A0(\pcpi_mul.rd[22] ),
    .A1(\pcpi_mul.rd[54] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _30041_ (.A0(_01908_),
    .A1(_01971_),
    .S(net481),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _30042_ (.A0(_01966_),
    .A1(_01965_),
    .S(_01714_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_2 _30043_ (.A0(_01968_),
    .A1(_01967_),
    .S(_01717_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_2 _30044_ (.A0(\pcpi_mul.rd[21] ),
    .A1(\pcpi_mul.rd[53] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _30045_ (.A0(_01908_),
    .A1(_01962_),
    .S(net481),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _30046_ (.A0(_01957_),
    .A1(_01956_),
    .S(net487),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_2 _30047_ (.A0(_01959_),
    .A1(_01958_),
    .S(_01717_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_2 _30048_ (.A0(\pcpi_mul.rd[20] ),
    .A1(\pcpi_mul.rd[52] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _30049_ (.A0(_01908_),
    .A1(_01953_),
    .S(net481),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _30050_ (.A0(_01948_),
    .A1(_01947_),
    .S(net487),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_2 _30051_ (.A0(_01950_),
    .A1(_01949_),
    .S(_01717_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_2 _30052_ (.A0(\pcpi_mul.rd[19] ),
    .A1(\pcpi_mul.rd[51] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_2 _30053_ (.A0(_01908_),
    .A1(_01944_),
    .S(net481),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _30054_ (.A0(_01939_),
    .A1(_01938_),
    .S(net487),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_2 _30055_ (.A0(_01941_),
    .A1(_01940_),
    .S(net446),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_2 _30056_ (.A0(\pcpi_mul.rd[18] ),
    .A1(\pcpi_mul.rd[50] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _30057_ (.A0(_01908_),
    .A1(_01935_),
    .S(net481),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_2 _30058_ (.A0(_01930_),
    .A1(_01929_),
    .S(net487),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_2 _30059_ (.A0(_01932_),
    .A1(_01931_),
    .S(net446),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_4 _30060_ (.A0(\pcpi_mul.rd[17] ),
    .A1(\pcpi_mul.rd[49] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_2 _30061_ (.A0(_01908_),
    .A1(_01926_),
    .S(net481),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _30062_ (.A0(_01921_),
    .A1(_01920_),
    .S(net487),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_2 _30063_ (.A0(_01923_),
    .A1(_01922_),
    .S(net446),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_2 _30064_ (.A0(\pcpi_mul.rd[16] ),
    .A1(\pcpi_mul.rd[48] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _30065_ (.A0(_01908_),
    .A1(_01917_),
    .S(net481),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _30066_ (.A0(_01912_),
    .A1(_01911_),
    .S(net487),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_2 _30067_ (.A0(_01914_),
    .A1(_01913_),
    .S(net446),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_2 _30068_ (.A0(\pcpi_mul.rd[15] ),
    .A1(\pcpi_mul.rd[47] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _30069_ (.A0(_01908_),
    .A1(_01907_),
    .S(_01816_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _30070_ (.A0(_01906_),
    .A1(_01904_),
    .S(net453),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _30071_ (.A0(net500),
    .A1(net57),
    .S(net317),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _30072_ (.A0(_01899_),
    .A1(_01898_),
    .S(net487),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_2 _30073_ (.A0(_01901_),
    .A1(_01900_),
    .S(_01717_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _30074_ (.A0(\pcpi_mul.rd[14] ),
    .A1(\pcpi_mul.rd[46] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_2 _30075_ (.A0(_01895_),
    .A1(_01894_),
    .S(_01816_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _30076_ (.A0(_01893_),
    .A1(_01891_),
    .S(net453),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _30077_ (.A0(net38),
    .A1(net497),
    .S(net317),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _30078_ (.A0(_01886_),
    .A1(_01885_),
    .S(net487),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_2 _30079_ (.A0(_01888_),
    .A1(_01887_),
    .S(net446),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_2 _30080_ (.A0(\pcpi_mul.rd[13] ),
    .A1(\pcpi_mul.rd[45] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _30081_ (.A0(_01882_),
    .A1(_01881_),
    .S(net481),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _30082_ (.A0(_01880_),
    .A1(_01878_),
    .S(net453),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _30083_ (.A0(net37),
    .A1(net54),
    .S(net317),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _30084_ (.A0(_01873_),
    .A1(_01872_),
    .S(net486),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_2 _30085_ (.A0(_01875_),
    .A1(_01874_),
    .S(net446),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _30086_ (.A0(\pcpi_mul.rd[12] ),
    .A1(\pcpi_mul.rd[44] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _30087_ (.A0(_01869_),
    .A1(_01868_),
    .S(net481),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _30088_ (.A0(_01867_),
    .A1(_01865_),
    .S(net453),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _30089_ (.A0(net36),
    .A1(net53),
    .S(net317),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _30090_ (.A0(_01860_),
    .A1(_01859_),
    .S(net486),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_2 _30091_ (.A0(_01862_),
    .A1(_01861_),
    .S(_01717_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_2 _30092_ (.A0(\pcpi_mul.rd[11] ),
    .A1(\pcpi_mul.rd[43] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_2 _30093_ (.A0(_01856_),
    .A1(_01855_),
    .S(net481),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _30094_ (.A0(_01854_),
    .A1(_01852_),
    .S(net453),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _30095_ (.A0(net35),
    .A1(net52),
    .S(net317),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _30096_ (.A0(_01847_),
    .A1(_01846_),
    .S(net486),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_2 _30097_ (.A0(_01849_),
    .A1(_01848_),
    .S(net446),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _30098_ (.A0(\pcpi_mul.rd[10] ),
    .A1(\pcpi_mul.rd[42] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _30099_ (.A0(_01843_),
    .A1(_01842_),
    .S(net481),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _30100_ (.A0(_01841_),
    .A1(_01839_),
    .S(net453),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _30101_ (.A0(net34),
    .A1(net51),
    .S(net317),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _30102_ (.A0(_01834_),
    .A1(_01833_),
    .S(net486),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_2 _30103_ (.A0(_01836_),
    .A1(_01835_),
    .S(net446),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_4 _30104_ (.A0(\pcpi_mul.rd[9] ),
    .A1(\pcpi_mul.rd[41] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_2 _30105_ (.A0(_01830_),
    .A1(_01829_),
    .S(net481),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _30106_ (.A0(_01828_),
    .A1(_01826_),
    .S(net453),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _30107_ (.A0(net64),
    .A1(net50),
    .S(net317),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _30108_ (.A0(_01821_),
    .A1(_01820_),
    .S(net486),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_2 _30109_ (.A0(_01823_),
    .A1(_01822_),
    .S(net446),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_2 _30110_ (.A0(\pcpi_mul.rd[8] ),
    .A1(\pcpi_mul.rd[40] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_2 _30111_ (.A0(_01817_),
    .A1(_01815_),
    .S(net481),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _30112_ (.A0(_01814_),
    .A1(_01812_),
    .S(net453),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _30113_ (.A0(net63),
    .A1(net49),
    .S(net317),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _30114_ (.A0(_01807_),
    .A1(_01806_),
    .S(net486),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_2 _30115_ (.A0(_01809_),
    .A1(_01808_),
    .S(net446),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_2 _30116_ (.A0(\pcpi_mul.rd[7] ),
    .A1(\pcpi_mul.rd[39] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _30117_ (.A0(_01803_),
    .A1(_01799_),
    .S(net453),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _30118_ (.A0(net62),
    .A1(net48),
    .S(net317),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _30119_ (.A0(_01800_),
    .A1(_01799_),
    .S(_00304_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _30120_ (.A0(_01794_),
    .A1(_01793_),
    .S(net485),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_2 _30121_ (.A0(_01796_),
    .A1(_01795_),
    .S(net446),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_2 _30122_ (.A0(\pcpi_mul.rd[6] ),
    .A1(\pcpi_mul.rd[38] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _30123_ (.A0(_01790_),
    .A1(_01786_),
    .S(net453),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _30124_ (.A0(net61),
    .A1(net47),
    .S(net317),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _30125_ (.A0(_01787_),
    .A1(_01786_),
    .S(_00304_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _30126_ (.A0(_01781_),
    .A1(_01780_),
    .S(net486),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_2 _30127_ (.A0(_01783_),
    .A1(_01782_),
    .S(net446),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_4 _30128_ (.A0(\pcpi_mul.rd[5] ),
    .A1(\pcpi_mul.rd[37] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_2 _30129_ (.A0(_01777_),
    .A1(_01773_),
    .S(net453),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _30130_ (.A0(net60),
    .A1(net46),
    .S(net317),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _30131_ (.A0(_01774_),
    .A1(_01773_),
    .S(_00304_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _30132_ (.A0(_01768_),
    .A1(_01767_),
    .S(net486),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_2 _30133_ (.A0(_01770_),
    .A1(_01769_),
    .S(net446),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_2 _30134_ (.A0(\pcpi_mul.rd[4] ),
    .A1(\pcpi_mul.rd[36] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_2 _30135_ (.A0(_01764_),
    .A1(_01760_),
    .S(net452),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _30136_ (.A0(net59),
    .A1(net45),
    .S(net317),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _30137_ (.A0(_01761_),
    .A1(_01760_),
    .S(_00304_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _30138_ (.A0(_01755_),
    .A1(_01754_),
    .S(net486),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_2 _30139_ (.A0(_01757_),
    .A1(_01756_),
    .S(net446),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_2 _30140_ (.A0(\pcpi_mul.rd[3] ),
    .A1(\pcpi_mul.rd[35] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_2 _30141_ (.A0(_01751_),
    .A1(_01747_),
    .S(net453),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _30142_ (.A0(net58),
    .A1(net498),
    .S(net317),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _30143_ (.A0(_01748_),
    .A1(_01747_),
    .S(_00304_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _30144_ (.A0(_01742_),
    .A1(_01741_),
    .S(net485),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_2 _30145_ (.A0(_01744_),
    .A1(_01743_),
    .S(net446),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_2 _30146_ (.A0(\pcpi_mul.rd[2] ),
    .A1(\pcpi_mul.rd[34] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_2 _30147_ (.A0(_01738_),
    .A1(_01734_),
    .S(net453),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _30148_ (.A0(net55),
    .A1(net42),
    .S(net317),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _30149_ (.A0(_01735_),
    .A1(_01734_),
    .S(_00304_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _30150_ (.A0(_01729_),
    .A1(_01728_),
    .S(net485),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _30151_ (.A0(_01731_),
    .A1(_01730_),
    .S(net446),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_2 _30152_ (.A0(\pcpi_mul.rd[1] ),
    .A1(\pcpi_mul.rd[33] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _30153_ (.A0(_01725_),
    .A1(_01721_),
    .S(net453),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _30154_ (.A0(net44),
    .A1(net499),
    .S(net317),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _30155_ (.A0(_01722_),
    .A1(_01721_),
    .S(_00304_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _30156_ (.A0(_01715_),
    .A1(_02559_),
    .S(net485),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_2 _30157_ (.A0(_01718_),
    .A1(_01716_),
    .S(net446),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_2 _30158_ (.A0(\pcpi_mul.rd[0] ),
    .A1(\pcpi_mul.rd[32] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_2 _30159_ (.A0(_01711_),
    .A1(_01707_),
    .S(net453),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _30160_ (.A0(net33),
    .A1(net40),
    .S(net317),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _30161_ (.A0(_01708_),
    .A1(_01707_),
    .S(_00304_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _30162_ (.A0(_01701_),
    .A1(_01696_),
    .S(_00311_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _30163_ (.A0(_01702_),
    .A1(_01696_),
    .S(\pcpi_mul.active[1] ),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _30164_ (.A0(_01696_),
    .A1(_01703_),
    .S(_00310_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _30165_ (.A0(_01693_),
    .A1(net273),
    .S(_00316_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _30166_ (.A0(_01690_),
    .A1(net272),
    .S(_00316_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _30167_ (.A0(_01687_),
    .A1(net271),
    .S(_00316_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _30168_ (.A0(_01684_),
    .A1(net270),
    .S(_00316_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _30169_ (.A0(\reg_next_pc[31] ),
    .A1(_01554_),
    .S(latched_store),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _30170_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(latched_stalu),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _30171_ (.A0(\reg_next_pc[30] ),
    .A1(_01551_),
    .S(latched_store),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _30172_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(latched_stalu),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _30173_ (.A0(\reg_next_pc[29] ),
    .A1(_01548_),
    .S(latched_store),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_2 _30174_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(latched_stalu),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _30175_ (.A0(\reg_next_pc[28] ),
    .A1(_01545_),
    .S(latched_store),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _30176_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(latched_stalu),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _30177_ (.A0(\reg_next_pc[27] ),
    .A1(_01542_),
    .S(latched_store),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_2 _30178_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(latched_stalu),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _30179_ (.A0(\reg_next_pc[26] ),
    .A1(_01539_),
    .S(latched_store),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _30180_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(latched_stalu),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _30181_ (.A0(\reg_next_pc[25] ),
    .A1(_01536_),
    .S(latched_store),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _30182_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(latched_stalu),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _30183_ (.A0(\reg_next_pc[24] ),
    .A1(_01533_),
    .S(latched_store),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_2 _30184_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(latched_stalu),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _30185_ (.A0(\reg_next_pc[23] ),
    .A1(_01530_),
    .S(latched_store),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _30186_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(latched_stalu),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _30187_ (.A0(\reg_next_pc[22] ),
    .A1(_01527_),
    .S(latched_store),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _30188_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(latched_stalu),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _30189_ (.A0(\reg_next_pc[21] ),
    .A1(_01524_),
    .S(latched_store),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _30190_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(latched_stalu),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _30191_ (.A0(\reg_next_pc[20] ),
    .A1(_01521_),
    .S(latched_store),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _30192_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(latched_stalu),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _30193_ (.A0(\reg_next_pc[19] ),
    .A1(_01518_),
    .S(latched_store),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_2 _30194_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(latched_stalu),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _30195_ (.A0(\reg_next_pc[18] ),
    .A1(_01515_),
    .S(latched_store),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _30196_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(latched_stalu),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _30197_ (.A0(\reg_next_pc[17] ),
    .A1(_01512_),
    .S(latched_store),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _30198_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(latched_stalu),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _30199_ (.A0(\reg_next_pc[16] ),
    .A1(_01509_),
    .S(latched_store),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _30200_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(latched_stalu),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _30201_ (.A0(\reg_next_pc[15] ),
    .A1(_01506_),
    .S(latched_store),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _30202_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(latched_stalu),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _30203_ (.A0(\reg_next_pc[14] ),
    .A1(_01503_),
    .S(latched_store),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _30204_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(latched_stalu),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _30205_ (.A0(\reg_next_pc[13] ),
    .A1(_01500_),
    .S(latched_store),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_2 _30206_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(latched_stalu),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _30207_ (.A0(\reg_next_pc[12] ),
    .A1(_01497_),
    .S(latched_store),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _30208_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(latched_stalu),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _30209_ (.A0(\reg_next_pc[11] ),
    .A1(_01494_),
    .S(latched_store),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_2 _30210_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(latched_stalu),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _30211_ (.A0(\reg_next_pc[10] ),
    .A1(_01491_),
    .S(latched_store),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _30212_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(latched_stalu),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _30213_ (.A0(\reg_next_pc[9] ),
    .A1(_01488_),
    .S(latched_store),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _30214_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(latched_stalu),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _30215_ (.A0(\reg_next_pc[8] ),
    .A1(_01485_),
    .S(latched_store),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _30216_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(latched_stalu),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _30217_ (.A0(\reg_next_pc[7] ),
    .A1(_01482_),
    .S(latched_store),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_2 _30218_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(latched_stalu),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _30219_ (.A0(\reg_next_pc[6] ),
    .A1(_01479_),
    .S(latched_store),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _30220_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(latched_stalu),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _30221_ (.A0(\reg_next_pc[5] ),
    .A1(_01476_),
    .S(latched_store),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_2 _30222_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(latched_stalu),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_4 _30223_ (.A0(_01474_),
    .A1(_01471_),
    .S(net455),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _30224_ (.A0(\reg_next_pc[4] ),
    .A1(_01472_),
    .S(latched_store),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _30225_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(latched_stalu),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _30226_ (.A0(\reg_next_pc[3] ),
    .A1(_01468_),
    .S(latched_store),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _30227_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _30228_ (.A0(\reg_next_pc[1] ),
    .A1(_01465_),
    .S(latched_store),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_2 _30229_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(latched_stalu),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _30230_ (.A0(_01301_),
    .A1(\timer[31] ),
    .S(_01208_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _30231_ (.A0(_01298_),
    .A1(\timer[30] ),
    .S(_01208_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _30232_ (.A0(_01295_),
    .A1(\timer[29] ),
    .S(_01208_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _30233_ (.A0(_01292_),
    .A1(\timer[28] ),
    .S(_01208_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _30234_ (.A0(_01289_),
    .A1(\timer[27] ),
    .S(net419),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _30235_ (.A0(_01286_),
    .A1(\timer[26] ),
    .S(net419),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _30236_ (.A0(_01283_),
    .A1(\timer[25] ),
    .S(net419),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _30237_ (.A0(_01280_),
    .A1(\timer[24] ),
    .S(net419),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _30238_ (.A0(_01277_),
    .A1(\timer[23] ),
    .S(net419),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _30239_ (.A0(_01274_),
    .A1(\timer[22] ),
    .S(net419),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _30240_ (.A0(_01271_),
    .A1(\timer[21] ),
    .S(net419),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _30241_ (.A0(_01268_),
    .A1(\timer[20] ),
    .S(net418),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _30242_ (.A0(_01265_),
    .A1(\timer[19] ),
    .S(net418),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _30243_ (.A0(_01262_),
    .A1(\timer[18] ),
    .S(net418),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _30244_ (.A0(_01259_),
    .A1(\timer[17] ),
    .S(net418),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _30245_ (.A0(_01256_),
    .A1(\timer[16] ),
    .S(net418),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _30246_ (.A0(_01253_),
    .A1(\timer[15] ),
    .S(net418),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _30247_ (.A0(_01250_),
    .A1(\timer[14] ),
    .S(net418),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _30248_ (.A0(_01247_),
    .A1(\timer[13] ),
    .S(net418),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _30249_ (.A0(_01244_),
    .A1(\timer[12] ),
    .S(net418),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _30250_ (.A0(_01241_),
    .A1(\timer[11] ),
    .S(net418),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _30251_ (.A0(_01238_),
    .A1(\timer[10] ),
    .S(net417),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _30252_ (.A0(_01235_),
    .A1(\timer[9] ),
    .S(net418),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _30253_ (.A0(_01232_),
    .A1(\timer[8] ),
    .S(net417),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _30254_ (.A0(_01229_),
    .A1(\timer[7] ),
    .S(net417),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _30255_ (.A0(_01226_),
    .A1(\timer[6] ),
    .S(net417),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _30256_ (.A0(_01223_),
    .A1(\timer[5] ),
    .S(net417),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _30257_ (.A0(_01220_),
    .A1(\timer[4] ),
    .S(net417),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _30258_ (.A0(_01217_),
    .A1(\timer[3] ),
    .S(net417),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _30259_ (.A0(_01214_),
    .A1(\timer[2] ),
    .S(net417),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _30260_ (.A0(_01211_),
    .A1(\timer[1] ),
    .S(net417),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_2 _30261_ (.A0(_01206_),
    .A1(_01201_),
    .S(net449),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_2 _30262_ (.A0(_01179_),
    .A1(_01174_),
    .S(net449),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_2 _30263_ (.A0(_01152_),
    .A1(_01147_),
    .S(net449),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_2 _30264_ (.A0(_01125_),
    .A1(_01120_),
    .S(net449),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_2 _30265_ (.A0(_01098_),
    .A1(_01093_),
    .S(net449),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_2 _30266_ (.A0(_01071_),
    .A1(_01066_),
    .S(net449),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_2 _30267_ (.A0(_01044_),
    .A1(_01039_),
    .S(net449),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_2 _30268_ (.A0(_01017_),
    .A1(_01012_),
    .S(net449),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_4 _30269_ (.A0(_00990_),
    .A1(_00985_),
    .S(net449),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_2 _30270_ (.A0(_00963_),
    .A1(_00958_),
    .S(net449),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_2 _30271_ (.A0(_00936_),
    .A1(_00931_),
    .S(net449),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_2 _30272_ (.A0(_00909_),
    .A1(_00904_),
    .S(net449),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_4 _30273_ (.A0(_00882_),
    .A1(_00877_),
    .S(net448),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_4 _30274_ (.A0(_00855_),
    .A1(_00850_),
    .S(net448),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_4 _30275_ (.A0(_00828_),
    .A1(_00823_),
    .S(net448),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_4 _30276_ (.A0(_00801_),
    .A1(_00796_),
    .S(net447),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_4 _30277_ (.A0(_00774_),
    .A1(_00769_),
    .S(net447),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_4 _30278_ (.A0(_00747_),
    .A1(_00742_),
    .S(net448),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_4 _30279_ (.A0(_00720_),
    .A1(_00715_),
    .S(net447),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_4 _30280_ (.A0(_00693_),
    .A1(_00688_),
    .S(net447),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_4 _30281_ (.A0(_00666_),
    .A1(_00661_),
    .S(net447),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_4 _30282_ (.A0(_00639_),
    .A1(_00634_),
    .S(net447),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_4 _30283_ (.A0(_00612_),
    .A1(_00607_),
    .S(net447),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_4 _30284_ (.A0(_00585_),
    .A1(_00580_),
    .S(net447),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_4 _30285_ (.A0(_00558_),
    .A1(_00553_),
    .S(net448),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_2 _30286_ (.A0(_00531_),
    .A1(_00526_),
    .S(net448),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_4 _30287_ (.A0(_00504_),
    .A1(_00499_),
    .S(net448),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_4 _30288_ (.A0(_00477_),
    .A1(_00472_),
    .S(net448),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_4 _30289_ (.A0(_00450_),
    .A1(_00445_),
    .S(net448),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_4 _30290_ (.A0(_00423_),
    .A1(_00418_),
    .S(net448),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_4 _30291_ (.A0(_00396_),
    .A1(_00391_),
    .S(net447),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_4 _30292_ (.A0(_00369_),
    .A1(_00365_),
    .S(net449),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_2 _30293_ (.A0(_00366_),
    .A1(_00367_),
    .S(net495),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_8 _30294_ (.A0(\decoded_rs1[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(net495),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_4 _30295_ (.A0(\decoded_rs1[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(net495),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_4 _30296_ (.A0(\decoded_rs1[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(net495),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_8 _30297_ (.A0(\decoded_rs1[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(net495),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _30298_ (.A0(_00349_),
    .A1(_00323_),
    .S(decoder_trigger),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _30299_ (.A0(_00350_),
    .A1(_00351_),
    .S(_00309_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _30300_ (.A0(_00352_),
    .A1(_00349_),
    .S(_00308_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _30301_ (.A0(_00355_),
    .A1(_00353_),
    .S(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _30302_ (.A0(_00337_),
    .A1(_00344_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _30303_ (.A0(_00345_),
    .A1(_00337_),
    .S(alu_wait),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_8 _30304_ (.A0(_00342_),
    .A1(_00340_),
    .S(_00341_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _30305_ (.A0(_00338_),
    .A1(_00337_),
    .S(_00296_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _30306_ (.A0(\mem_rdata_q[12] ),
    .A1(_00334_),
    .S(\mem_rdata_q[13] ),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _30307_ (.A0(\cpu_state[1] ),
    .A1(_00302_),
    .S(\cpu_state[4] ),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _30308_ (.A0(_00322_),
    .A1(_00296_),
    .S(\cpu_state[6] ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_2 _30309_ (.A0(_00315_),
    .A1(alu_wait),
    .S(\cpu_state[4] ),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_2 _30310_ (.A0(\mem_rdata_q[6] ),
    .A1(net61),
    .S(net445),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_4 _30311_ (.A0(\mem_rdata_q[5] ),
    .A1(net60),
    .S(net445),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_2 _30312_ (.A0(\mem_rdata_q[4] ),
    .A1(net59),
    .S(net445),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _30313_ (.A0(\mem_rdata_q[3] ),
    .A1(net58),
    .S(mem_xfer),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _30314_ (.A0(\mem_rdata_q[2] ),
    .A1(net55),
    .S(net445),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_2 _30315_ (.A0(\mem_rdata_q[1] ),
    .A1(net44),
    .S(net445),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_2 _30316_ (.A0(\mem_rdata_q[0] ),
    .A1(net33),
    .S(mem_xfer),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _30317_ (.A0(\cpu_state[1] ),
    .A1(instr_retirq),
    .S(\cpu_state[2] ),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _30318_ (.A0(_00319_),
    .A1(\cpu_state[5] ),
    .S(_00296_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _30319_ (.A0(_00317_),
    .A1(\cpu_state[6] ),
    .S(_00296_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _30320_ (.A0(_00313_),
    .A1(_00312_),
    .S(_00307_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _30321_ (.A0(_00298_),
    .A1(_00299_),
    .S(_00289_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _30322_ (.A0(\reg_next_pc[2] ),
    .A1(_00293_),
    .S(latched_store),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _30323_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _30324_ (.A0(_00126_),
    .A1(_00122_),
    .S(net489),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _30325_ (.A0(_00120_),
    .A1(_00116_),
    .S(net489),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _30326_ (.A0(_00114_),
    .A1(_00110_),
    .S(net489),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _30327_ (.A0(_00108_),
    .A1(_00104_),
    .S(net225),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _30328_ (.A0(_00102_),
    .A1(_00095_),
    .S(net489),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _30329_ (.A0(_00092_),
    .A1(_00085_),
    .S(net489),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _30330_ (.A0(_00082_),
    .A1(_00068_),
    .S(net489),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _30331_ (.A0(_00064_),
    .A1(_00050_),
    .S(net489),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _30332_ (.A0(_01694_),
    .A1(_01695_),
    .S(_00290_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _30333_ (.A0(_01691_),
    .A1(_01692_),
    .S(_00290_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _30334_ (.A0(_01688_),
    .A1(_01689_),
    .S(_00290_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _30335_ (.A0(_01685_),
    .A1(_01686_),
    .S(_00290_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _30336_ (.A0(_01679_),
    .A1(_01680_),
    .S(instr_jal),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _30337_ (.A0(_01682_),
    .A1(_02581_),
    .S(net416),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _30338_ (.A0(_01675_),
    .A1(_01676_),
    .S(instr_jal),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _30339_ (.A0(_01678_),
    .A1(_02580_),
    .S(net416),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _30340_ (.A0(_01671_),
    .A1(_01672_),
    .S(instr_jal),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _30341_ (.A0(_01674_),
    .A1(_02579_),
    .S(net416),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _30342_ (.A0(_01667_),
    .A1(_01668_),
    .S(instr_jal),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _30343_ (.A0(_01670_),
    .A1(_02578_),
    .S(net416),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _30344_ (.A0(_01663_),
    .A1(_01664_),
    .S(instr_jal),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _30345_ (.A0(_01666_),
    .A1(_02577_),
    .S(net416),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _30346_ (.A0(_01659_),
    .A1(_01660_),
    .S(instr_jal),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _30347_ (.A0(_01662_),
    .A1(_02576_),
    .S(net416),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _30348_ (.A0(_01655_),
    .A1(_01656_),
    .S(instr_jal),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _30349_ (.A0(_01658_),
    .A1(_02575_),
    .S(net416),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _30350_ (.A0(_01651_),
    .A1(_01652_),
    .S(instr_jal),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _30351_ (.A0(_01654_),
    .A1(_02574_),
    .S(net416),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _30352_ (.A0(_01647_),
    .A1(_01648_),
    .S(instr_jal),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _30353_ (.A0(_01650_),
    .A1(_02573_),
    .S(net416),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _30354_ (.A0(_01643_),
    .A1(_01644_),
    .S(instr_jal),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _30355_ (.A0(_01646_),
    .A1(_02572_),
    .S(net416),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _30356_ (.A0(_01639_),
    .A1(_01640_),
    .S(instr_jal),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _30357_ (.A0(_01642_),
    .A1(_02570_),
    .S(net416),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _30358_ (.A0(_01635_),
    .A1(_01636_),
    .S(instr_jal),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _30359_ (.A0(_01638_),
    .A1(_02569_),
    .S(net416),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _30360_ (.A0(_01631_),
    .A1(_01632_),
    .S(instr_jal),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _30361_ (.A0(_01634_),
    .A1(_02568_),
    .S(net416),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _30362_ (.A0(_01627_),
    .A1(_01628_),
    .S(instr_jal),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _30363_ (.A0(_01630_),
    .A1(_02567_),
    .S(net416),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _30364_ (.A0(_01623_),
    .A1(_01624_),
    .S(instr_jal),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _30365_ (.A0(_01626_),
    .A1(_02566_),
    .S(net416),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _30366_ (.A0(_01619_),
    .A1(_01620_),
    .S(instr_jal),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _30367_ (.A0(_01622_),
    .A1(_02565_),
    .S(net416),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _30368_ (.A0(_01615_),
    .A1(_01616_),
    .S(instr_jal),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _30369_ (.A0(_01618_),
    .A1(_02564_),
    .S(net416),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _30370_ (.A0(_01611_),
    .A1(_01612_),
    .S(instr_jal),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _30371_ (.A0(_01614_),
    .A1(_02563_),
    .S(net416),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _30372_ (.A0(_01607_),
    .A1(_01608_),
    .S(instr_jal),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _30373_ (.A0(_01610_),
    .A1(_02562_),
    .S(net416),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _30374_ (.A0(_01603_),
    .A1(_01604_),
    .S(instr_jal),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _30375_ (.A0(_01606_),
    .A1(_02561_),
    .S(_00308_),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _30376_ (.A0(_01599_),
    .A1(_01600_),
    .S(instr_jal),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _30377_ (.A0(_01602_),
    .A1(_02589_),
    .S(_00308_),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _30378_ (.A0(_01595_),
    .A1(_01596_),
    .S(instr_jal),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _30379_ (.A0(_01598_),
    .A1(_02588_),
    .S(_00308_),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _30380_ (.A0(_01591_),
    .A1(_01592_),
    .S(instr_jal),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _30381_ (.A0(_01594_),
    .A1(_02587_),
    .S(net416),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _30382_ (.A0(_01587_),
    .A1(_01588_),
    .S(instr_jal),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _30383_ (.A0(_01590_),
    .A1(_02586_),
    .S(_00308_),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _30384_ (.A0(_01583_),
    .A1(_01584_),
    .S(instr_jal),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _30385_ (.A0(_01586_),
    .A1(_02585_),
    .S(_00308_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _30386_ (.A0(_01579_),
    .A1(_01580_),
    .S(instr_jal),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _30387_ (.A0(_01582_),
    .A1(_02584_),
    .S(_00308_),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _30388_ (.A0(_01575_),
    .A1(_01576_),
    .S(instr_jal),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _30389_ (.A0(_01578_),
    .A1(_02583_),
    .S(_00308_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _30390_ (.A0(_01571_),
    .A1(_01572_),
    .S(instr_jal),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _30391_ (.A0(_01574_),
    .A1(_02582_),
    .S(_00308_),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _30392_ (.A0(_01567_),
    .A1(_01568_),
    .S(instr_jal),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _30393_ (.A0(_01570_),
    .A1(_02571_),
    .S(_00308_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _30394_ (.A0(_01561_),
    .A1(_01562_),
    .S(instr_jal),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _30395_ (.A0(_02560_),
    .A1(_01563_),
    .S(decoder_trigger),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _30396_ (.A0(_01564_),
    .A1(_01565_),
    .S(_00309_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _30397_ (.A0(_01566_),
    .A1(_02560_),
    .S(_00308_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _30398_ (.A0(_02590_),
    .A1(_01557_),
    .S(instr_jal),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _30399_ (.A0(_02590_),
    .A1(_01558_),
    .S(decoder_trigger),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _30400_ (.A0(_01559_),
    .A1(_02590_),
    .S(_00309_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _30401_ (.A0(_01560_),
    .A1(_02590_),
    .S(_00308_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _30402_ (.A0(\cpuregs_rs1[31] ),
    .A1(_01462_),
    .S(is_lui_auipc_jal),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _30403_ (.A0(_01464_),
    .A1(_01463_),
    .S(net484),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _30404_ (.A0(\cpuregs_rs1[30] ),
    .A1(_01459_),
    .S(is_lui_auipc_jal),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _30405_ (.A0(_01461_),
    .A1(_01460_),
    .S(net484),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _30406_ (.A0(\cpuregs_rs1[29] ),
    .A1(_01456_),
    .S(is_lui_auipc_jal),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _30407_ (.A0(_01458_),
    .A1(_01457_),
    .S(net484),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _30408_ (.A0(\cpuregs_rs1[28] ),
    .A1(_01453_),
    .S(is_lui_auipc_jal),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _30409_ (.A0(_01455_),
    .A1(_01454_),
    .S(net484),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _30410_ (.A0(\cpuregs_rs1[27] ),
    .A1(_01450_),
    .S(is_lui_auipc_jal),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _30411_ (.A0(_01452_),
    .A1(_01451_),
    .S(net484),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _30412_ (.A0(\cpuregs_rs1[26] ),
    .A1(_01447_),
    .S(is_lui_auipc_jal),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _30413_ (.A0(_01449_),
    .A1(_01448_),
    .S(net484),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _30414_ (.A0(\cpuregs_rs1[25] ),
    .A1(_01444_),
    .S(is_lui_auipc_jal),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _30415_ (.A0(_01446_),
    .A1(_01445_),
    .S(net484),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _30416_ (.A0(\cpuregs_rs1[24] ),
    .A1(_01441_),
    .S(is_lui_auipc_jal),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _30417_ (.A0(_01443_),
    .A1(_01442_),
    .S(net484),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _30418_ (.A0(\cpuregs_rs1[23] ),
    .A1(_01438_),
    .S(is_lui_auipc_jal),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _30419_ (.A0(_01440_),
    .A1(_01439_),
    .S(net484),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_2 _30420_ (.A0(\cpuregs_rs1[22] ),
    .A1(_01435_),
    .S(is_lui_auipc_jal),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _30421_ (.A0(_01437_),
    .A1(_01436_),
    .S(net484),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_2 _30422_ (.A0(\cpuregs_rs1[21] ),
    .A1(_01432_),
    .S(is_lui_auipc_jal),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _30423_ (.A0(_01434_),
    .A1(_01433_),
    .S(net484),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_2 _30424_ (.A0(\cpuregs_rs1[20] ),
    .A1(_01429_),
    .S(is_lui_auipc_jal),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _30425_ (.A0(_01431_),
    .A1(_01430_),
    .S(net484),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _30426_ (.A0(\cpuregs_rs1[19] ),
    .A1(_01426_),
    .S(is_lui_auipc_jal),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _30427_ (.A0(_01428_),
    .A1(_01427_),
    .S(net483),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _30428_ (.A0(\cpuregs_rs1[18] ),
    .A1(_01423_),
    .S(is_lui_auipc_jal),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _30429_ (.A0(_01425_),
    .A1(_01424_),
    .S(net483),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _30430_ (.A0(\cpuregs_rs1[17] ),
    .A1(_01420_),
    .S(is_lui_auipc_jal),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _30431_ (.A0(_01422_),
    .A1(_01421_),
    .S(net483),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _30432_ (.A0(\cpuregs_rs1[16] ),
    .A1(_01417_),
    .S(is_lui_auipc_jal),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _30433_ (.A0(_01419_),
    .A1(_01418_),
    .S(net483),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _30434_ (.A0(\cpuregs_rs1[15] ),
    .A1(_01414_),
    .S(is_lui_auipc_jal),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _30435_ (.A0(_01416_),
    .A1(_01415_),
    .S(net483),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _30436_ (.A0(\cpuregs_rs1[14] ),
    .A1(_01411_),
    .S(is_lui_auipc_jal),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _30437_ (.A0(_01413_),
    .A1(_01412_),
    .S(net483),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _30438_ (.A0(\cpuregs_rs1[13] ),
    .A1(_01408_),
    .S(is_lui_auipc_jal),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _30439_ (.A0(_01410_),
    .A1(_01409_),
    .S(net483),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _30440_ (.A0(\cpuregs_rs1[12] ),
    .A1(_01405_),
    .S(is_lui_auipc_jal),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _30441_ (.A0(_01407_),
    .A1(_01406_),
    .S(net483),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _30442_ (.A0(\cpuregs_rs1[11] ),
    .A1(_01402_),
    .S(is_lui_auipc_jal),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _30443_ (.A0(_01404_),
    .A1(_01403_),
    .S(net483),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _30444_ (.A0(\cpuregs_rs1[10] ),
    .A1(_01399_),
    .S(is_lui_auipc_jal),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _30445_ (.A0(_01401_),
    .A1(_01400_),
    .S(net483),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _30446_ (.A0(\cpuregs_rs1[9] ),
    .A1(_01396_),
    .S(is_lui_auipc_jal),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _30447_ (.A0(_01398_),
    .A1(_01397_),
    .S(net483),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _30448_ (.A0(\cpuregs_rs1[8] ),
    .A1(_01393_),
    .S(is_lui_auipc_jal),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _30449_ (.A0(_01395_),
    .A1(_01394_),
    .S(net483),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _30450_ (.A0(\cpuregs_rs1[7] ),
    .A1(_01390_),
    .S(is_lui_auipc_jal),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _30451_ (.A0(_01392_),
    .A1(_01391_),
    .S(net483),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _30452_ (.A0(\cpuregs_rs1[6] ),
    .A1(_01387_),
    .S(is_lui_auipc_jal),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _30453_ (.A0(_01389_),
    .A1(_01388_),
    .S(net483),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _30454_ (.A0(\cpuregs_rs1[5] ),
    .A1(_01384_),
    .S(is_lui_auipc_jal),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _30455_ (.A0(_01386_),
    .A1(_01385_),
    .S(net483),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _30456_ (.A0(\cpuregs_rs1[4] ),
    .A1(_01381_),
    .S(is_lui_auipc_jal),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _30457_ (.A0(_01383_),
    .A1(_01382_),
    .S(net483),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _30458_ (.A0(\cpuregs_rs1[3] ),
    .A1(_01378_),
    .S(is_lui_auipc_jal),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _30459_ (.A0(_01380_),
    .A1(_01379_),
    .S(net484),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _30460_ (.A0(\cpuregs_rs1[2] ),
    .A1(_01375_),
    .S(is_lui_auipc_jal),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _30461_ (.A0(_01377_),
    .A1(_01376_),
    .S(net484),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _30462_ (.A0(\cpuregs_rs1[1] ),
    .A1(_01372_),
    .S(is_lui_auipc_jal),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _30463_ (.A0(_01374_),
    .A1(_01373_),
    .S(_00297_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _30464_ (.A0(\cpuregs_rs1[0] ),
    .A1(_01369_),
    .S(is_lui_auipc_jal),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _30465_ (.A0(_01371_),
    .A1(_01370_),
    .S(_00297_),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _30466_ (.A0(_01367_),
    .A1(\decoded_imm[31] ),
    .S(_01304_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _30467_ (.A0(_01368_),
    .A1(\cpuregs_rs1[31] ),
    .S(net495),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _30468_ (.A0(_01365_),
    .A1(\decoded_imm[30] ),
    .S(_01304_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _30469_ (.A0(_01366_),
    .A1(\cpuregs_rs1[30] ),
    .S(net495),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _30470_ (.A0(_01363_),
    .A1(\decoded_imm[29] ),
    .S(_01304_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _30471_ (.A0(_01364_),
    .A1(\cpuregs_rs1[29] ),
    .S(net495),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _30472_ (.A0(_01361_),
    .A1(\decoded_imm[28] ),
    .S(_01304_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _30473_ (.A0(_01362_),
    .A1(\cpuregs_rs1[28] ),
    .S(net495),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _30474_ (.A0(_01359_),
    .A1(\decoded_imm[27] ),
    .S(_01304_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _30475_ (.A0(_01360_),
    .A1(\cpuregs_rs1[27] ),
    .S(net495),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _30476_ (.A0(_01357_),
    .A1(\decoded_imm[26] ),
    .S(_01304_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _30477_ (.A0(_01358_),
    .A1(\cpuregs_rs1[26] ),
    .S(net495),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _30478_ (.A0(_01355_),
    .A1(\decoded_imm[25] ),
    .S(_01304_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _30479_ (.A0(_01356_),
    .A1(\cpuregs_rs1[25] ),
    .S(net495),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _30480_ (.A0(_01353_),
    .A1(\decoded_imm[24] ),
    .S(_01304_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _30481_ (.A0(_01354_),
    .A1(\cpuregs_rs1[24] ),
    .S(net495),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _30482_ (.A0(_01351_),
    .A1(\decoded_imm[23] ),
    .S(net482),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _30483_ (.A0(_01352_),
    .A1(\cpuregs_rs1[23] ),
    .S(net495),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _30484_ (.A0(_01349_),
    .A1(\decoded_imm[22] ),
    .S(net482),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _30485_ (.A0(_01350_),
    .A1(\cpuregs_rs1[22] ),
    .S(net495),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _30486_ (.A0(_01347_),
    .A1(\decoded_imm[21] ),
    .S(net482),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _30487_ (.A0(_01348_),
    .A1(\cpuregs_rs1[21] ),
    .S(net495),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _30488_ (.A0(_01345_),
    .A1(\decoded_imm[20] ),
    .S(net482),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _30489_ (.A0(_01346_),
    .A1(\cpuregs_rs1[20] ),
    .S(net495),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _30490_ (.A0(_01343_),
    .A1(\decoded_imm[19] ),
    .S(net482),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _30491_ (.A0(_01344_),
    .A1(\cpuregs_rs1[19] ),
    .S(net495),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _30492_ (.A0(_01341_),
    .A1(\decoded_imm[18] ),
    .S(net482),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _30493_ (.A0(_01342_),
    .A1(\cpuregs_rs1[18] ),
    .S(net495),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _30494_ (.A0(_01339_),
    .A1(\decoded_imm[17] ),
    .S(net482),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _30495_ (.A0(_01340_),
    .A1(\cpuregs_rs1[17] ),
    .S(net495),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _30496_ (.A0(_01337_),
    .A1(\decoded_imm[16] ),
    .S(net482),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _30497_ (.A0(_01338_),
    .A1(\cpuregs_rs1[16] ),
    .S(net495),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _30498_ (.A0(_01335_),
    .A1(\decoded_imm[15] ),
    .S(net482),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _30499_ (.A0(_01336_),
    .A1(\cpuregs_rs1[15] ),
    .S(net495),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _30500_ (.A0(_01333_),
    .A1(\decoded_imm[14] ),
    .S(net482),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _30501_ (.A0(_01334_),
    .A1(\cpuregs_rs1[14] ),
    .S(net495),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _30502_ (.A0(_01331_),
    .A1(\decoded_imm[13] ),
    .S(net482),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _30503_ (.A0(_01332_),
    .A1(\cpuregs_rs1[13] ),
    .S(net495),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _30504_ (.A0(_01329_),
    .A1(\decoded_imm[12] ),
    .S(net482),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _30505_ (.A0(_01330_),
    .A1(\cpuregs_rs1[12] ),
    .S(net495),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _30506_ (.A0(_01327_),
    .A1(\decoded_imm[11] ),
    .S(net482),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _30507_ (.A0(_01328_),
    .A1(\cpuregs_rs1[11] ),
    .S(net495),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _30508_ (.A0(_01325_),
    .A1(\decoded_imm[10] ),
    .S(net482),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _30509_ (.A0(_01326_),
    .A1(\cpuregs_rs1[10] ),
    .S(net495),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _30510_ (.A0(_01323_),
    .A1(\decoded_imm[9] ),
    .S(net482),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _30511_ (.A0(_01324_),
    .A1(\cpuregs_rs1[9] ),
    .S(net495),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _30512_ (.A0(_01321_),
    .A1(\decoded_imm[8] ),
    .S(net482),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _30513_ (.A0(_01322_),
    .A1(\cpuregs_rs1[8] ),
    .S(net495),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _30514_ (.A0(_01319_),
    .A1(\decoded_imm[7] ),
    .S(net482),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _30515_ (.A0(_01320_),
    .A1(\cpuregs_rs1[7] ),
    .S(net495),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _30516_ (.A0(_01317_),
    .A1(\decoded_imm[6] ),
    .S(net482),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _30517_ (.A0(_01318_),
    .A1(\cpuregs_rs1[6] ),
    .S(net495),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _30518_ (.A0(_01315_),
    .A1(\decoded_imm[5] ),
    .S(net482),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _30519_ (.A0(_01316_),
    .A1(\cpuregs_rs1[5] ),
    .S(net495),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _30520_ (.A0(\decoded_imm[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(is_slli_srli_srai),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _30521_ (.A0(_01313_),
    .A1(\decoded_imm[4] ),
    .S(_01304_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _30522_ (.A0(_01314_),
    .A1(\cpuregs_rs1[4] ),
    .S(net495),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _30523_ (.A0(\decoded_imm[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(is_slli_srli_srai),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _30524_ (.A0(_01311_),
    .A1(\decoded_imm[3] ),
    .S(_01304_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _30525_ (.A0(_01312_),
    .A1(\cpuregs_rs1[3] ),
    .S(net495),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _30526_ (.A0(\decoded_imm[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(is_slli_srli_srai),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _30527_ (.A0(_01309_),
    .A1(\decoded_imm[2] ),
    .S(_01304_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _30528_ (.A0(_01310_),
    .A1(\cpuregs_rs1[2] ),
    .S(net495),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _30529_ (.A0(\decoded_imm[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(is_slli_srli_srai),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _30530_ (.A0(_01307_),
    .A1(\decoded_imm[1] ),
    .S(_01304_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _30531_ (.A0(_01308_),
    .A1(\cpuregs_rs1[1] ),
    .S(net495),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _30532_ (.A0(\decoded_imm[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(is_slli_srli_srai),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _30533_ (.A0(_01305_),
    .A1(\decoded_imm[0] ),
    .S(_01304_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _30534_ (.A0(_01306_),
    .A1(\cpuregs_rs1[0] ),
    .S(net495),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _30535_ (.A0(_01302_),
    .A1(\cpuregs_rs1[31] ),
    .S(net494),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _30536_ (.A0(_01302_),
    .A1(_01303_),
    .S(\cpu_state[2] ),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _30537_ (.A0(_01299_),
    .A1(\cpuregs_rs1[30] ),
    .S(net494),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _30538_ (.A0(_01299_),
    .A1(_01300_),
    .S(\cpu_state[2] ),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _30539_ (.A0(_01296_),
    .A1(\cpuregs_rs1[29] ),
    .S(net494),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _30540_ (.A0(_01296_),
    .A1(_01297_),
    .S(\cpu_state[2] ),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _30541_ (.A0(_01293_),
    .A1(\cpuregs_rs1[28] ),
    .S(net494),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _30542_ (.A0(_01293_),
    .A1(_01294_),
    .S(\cpu_state[2] ),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _30543_ (.A0(_01290_),
    .A1(\cpuregs_rs1[27] ),
    .S(net494),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _30544_ (.A0(_01290_),
    .A1(_01291_),
    .S(\cpu_state[2] ),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _30545_ (.A0(_01287_),
    .A1(\cpuregs_rs1[26] ),
    .S(net494),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _30546_ (.A0(_01287_),
    .A1(_01288_),
    .S(\cpu_state[2] ),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _30547_ (.A0(_01284_),
    .A1(\cpuregs_rs1[25] ),
    .S(net494),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _30548_ (.A0(_01284_),
    .A1(_01285_),
    .S(\cpu_state[2] ),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _30549_ (.A0(_01281_),
    .A1(\cpuregs_rs1[24] ),
    .S(net494),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _30550_ (.A0(_01281_),
    .A1(_01282_),
    .S(\cpu_state[2] ),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _30551_ (.A0(_01278_),
    .A1(\cpuregs_rs1[23] ),
    .S(net494),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _30552_ (.A0(_01278_),
    .A1(_01279_),
    .S(\cpu_state[2] ),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _30553_ (.A0(_01275_),
    .A1(\cpuregs_rs1[22] ),
    .S(net494),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _30554_ (.A0(_01275_),
    .A1(_01276_),
    .S(\cpu_state[2] ),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _30555_ (.A0(_01272_),
    .A1(\cpuregs_rs1[21] ),
    .S(net494),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _30556_ (.A0(_01272_),
    .A1(_01273_),
    .S(\cpu_state[2] ),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _30557_ (.A0(_01269_),
    .A1(\cpuregs_rs1[20] ),
    .S(net494),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _30558_ (.A0(_01269_),
    .A1(_01270_),
    .S(\cpu_state[2] ),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _30559_ (.A0(_01266_),
    .A1(\cpuregs_rs1[19] ),
    .S(net494),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _30560_ (.A0(_01266_),
    .A1(_01267_),
    .S(\cpu_state[2] ),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _30561_ (.A0(_01263_),
    .A1(\cpuregs_rs1[18] ),
    .S(net494),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _30562_ (.A0(_01263_),
    .A1(_01264_),
    .S(\cpu_state[2] ),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _30563_ (.A0(_01260_),
    .A1(\cpuregs_rs1[17] ),
    .S(net494),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _30564_ (.A0(_01260_),
    .A1(_01261_),
    .S(\cpu_state[2] ),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _30565_ (.A0(_01257_),
    .A1(\cpuregs_rs1[16] ),
    .S(net494),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _30566_ (.A0(_01257_),
    .A1(_01258_),
    .S(\cpu_state[2] ),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _30567_ (.A0(_01254_),
    .A1(\cpuregs_rs1[15] ),
    .S(net494),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _30568_ (.A0(_01254_),
    .A1(_01255_),
    .S(\cpu_state[2] ),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _30569_ (.A0(_01251_),
    .A1(\cpuregs_rs1[14] ),
    .S(net494),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _30570_ (.A0(_01251_),
    .A1(_01252_),
    .S(\cpu_state[2] ),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _30571_ (.A0(_01248_),
    .A1(\cpuregs_rs1[13] ),
    .S(net494),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _30572_ (.A0(_01248_),
    .A1(_01249_),
    .S(\cpu_state[2] ),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _30573_ (.A0(_01245_),
    .A1(\cpuregs_rs1[12] ),
    .S(net494),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _30574_ (.A0(_01245_),
    .A1(_01246_),
    .S(\cpu_state[2] ),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _30575_ (.A0(_01242_),
    .A1(\cpuregs_rs1[11] ),
    .S(net494),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _30576_ (.A0(_01242_),
    .A1(_01243_),
    .S(\cpu_state[2] ),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _30577_ (.A0(_01239_),
    .A1(\cpuregs_rs1[10] ),
    .S(net494),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _30578_ (.A0(_01239_),
    .A1(_01240_),
    .S(\cpu_state[2] ),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _30579_ (.A0(_01236_),
    .A1(\cpuregs_rs1[9] ),
    .S(net494),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _30580_ (.A0(_01236_),
    .A1(_01237_),
    .S(\cpu_state[2] ),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _30581_ (.A0(_01233_),
    .A1(\cpuregs_rs1[8] ),
    .S(net494),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _30582_ (.A0(_01233_),
    .A1(_01234_),
    .S(\cpu_state[2] ),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _30583_ (.A0(_01230_),
    .A1(\cpuregs_rs1[7] ),
    .S(net494),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _30584_ (.A0(_01230_),
    .A1(_01231_),
    .S(\cpu_state[2] ),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _30585_ (.A0(_01227_),
    .A1(\cpuregs_rs1[6] ),
    .S(net494),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _30586_ (.A0(_01227_),
    .A1(_01228_),
    .S(\cpu_state[2] ),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _30587_ (.A0(_01224_),
    .A1(\cpuregs_rs1[5] ),
    .S(net494),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _30588_ (.A0(_01224_),
    .A1(_01225_),
    .S(\cpu_state[2] ),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _30589_ (.A0(_01221_),
    .A1(\cpuregs_rs1[4] ),
    .S(net494),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _30590_ (.A0(_01221_),
    .A1(_01222_),
    .S(\cpu_state[2] ),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _30591_ (.A0(_01218_),
    .A1(\cpuregs_rs1[3] ),
    .S(net494),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _30592_ (.A0(_01218_),
    .A1(_01219_),
    .S(\cpu_state[2] ),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _30593_ (.A0(_01215_),
    .A1(\cpuregs_rs1[2] ),
    .S(net494),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _30594_ (.A0(_01215_),
    .A1(_01216_),
    .S(\cpu_state[2] ),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _30595_ (.A0(_01212_),
    .A1(\cpuregs_rs1[1] ),
    .S(net494),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _30596_ (.A0(_01212_),
    .A1(_01213_),
    .S(\cpu_state[2] ),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _30597_ (.A0(_01209_),
    .A1(\cpuregs_rs1[0] ),
    .S(net494),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _30598_ (.A0(_01209_),
    .A1(_01210_),
    .S(\cpu_state[2] ),
    .X(_02411_));
 sky130_fd_sc_hd__mux4_1 _30599_ (.A0(_01202_),
    .A1(_01203_),
    .A2(_01204_),
    .A3(_01205_),
    .S0(net464),
    .S1(net472),
    .X(_01206_));
 sky130_fd_sc_hd__mux4_2 _30600_ (.A0(_01181_),
    .A1(_01182_),
    .A2(_01183_),
    .A3(_01184_),
    .S0(net465),
    .S1(net472),
    .X(_01185_));
 sky130_fd_sc_hd__mux4_2 _30601_ (.A0(_01186_),
    .A1(_01187_),
    .A2(_01188_),
    .A3(_01189_),
    .S0(net465),
    .S1(net472),
    .X(_01190_));
 sky130_fd_sc_hd__mux4_1 _30602_ (.A0(_01191_),
    .A1(_01192_),
    .A2(_01193_),
    .A3(_01194_),
    .S0(net465),
    .S1(net472),
    .X(_01195_));
 sky130_fd_sc_hd__mux4_1 _30603_ (.A0(_01196_),
    .A1(_01197_),
    .A2(_01198_),
    .A3(_01199_),
    .S0(net464),
    .S1(net472),
    .X(_01200_));
 sky130_fd_sc_hd__mux4_2 _30604_ (.A0(_01185_),
    .A1(_01190_),
    .A2(_01195_),
    .A3(_01200_),
    .S0(net477),
    .S1(net480),
    .X(_01201_));
 sky130_fd_sc_hd__mux4_1 _30605_ (.A0(_01175_),
    .A1(_01176_),
    .A2(_01177_),
    .A3(_01178_),
    .S0(net464),
    .S1(net472),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_2 _30606_ (.A0(_01154_),
    .A1(_01155_),
    .A2(_01156_),
    .A3(_01157_),
    .S0(net464),
    .S1(net472),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_2 _30607_ (.A0(_01159_),
    .A1(_01160_),
    .A2(_01161_),
    .A3(_01162_),
    .S0(net464),
    .S1(net472),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_2 _30608_ (.A0(_01164_),
    .A1(_01165_),
    .A2(_01166_),
    .A3(_01167_),
    .S0(net464),
    .S1(net472),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_1 _30609_ (.A0(_01169_),
    .A1(_01170_),
    .A2(_01171_),
    .A3(_01172_),
    .S0(net464),
    .S1(net472),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_2 _30610_ (.A0(_01158_),
    .A1(_01163_),
    .A2(_01168_),
    .A3(_01173_),
    .S0(net477),
    .S1(net480),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_1 _30611_ (.A0(_01148_),
    .A1(_01149_),
    .A2(_01150_),
    .A3(_01151_),
    .S0(net465),
    .S1(net472),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_1 _30612_ (.A0(_01127_),
    .A1(_01128_),
    .A2(_01129_),
    .A3(_01130_),
    .S0(net465),
    .S1(net473),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_1 _30613_ (.A0(_01132_),
    .A1(_01133_),
    .A2(_01134_),
    .A3(_01135_),
    .S0(net465),
    .S1(net473),
    .X(_01136_));
 sky130_fd_sc_hd__mux4_1 _30614_ (.A0(_01137_),
    .A1(_01138_),
    .A2(_01139_),
    .A3(_01140_),
    .S0(net465),
    .S1(net473),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_2 _30615_ (.A0(_01142_),
    .A1(_01143_),
    .A2(_01144_),
    .A3(_01145_),
    .S0(net465),
    .S1(net472),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_2 _30616_ (.A0(_01131_),
    .A1(_01136_),
    .A2(_01141_),
    .A3(_01146_),
    .S0(net477),
    .S1(net480),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_1 _30617_ (.A0(_01121_),
    .A1(_01122_),
    .A2(_01123_),
    .A3(_01124_),
    .S0(net465),
    .S1(net472),
    .X(_01125_));
 sky130_fd_sc_hd__mux4_1 _30618_ (.A0(_01100_),
    .A1(_01101_),
    .A2(_01102_),
    .A3(_01103_),
    .S0(net464),
    .S1(net472),
    .X(_01104_));
 sky130_fd_sc_hd__mux4_2 _30619_ (.A0(_01105_),
    .A1(_01106_),
    .A2(_01107_),
    .A3(_01108_),
    .S0(net464),
    .S1(net472),
    .X(_01109_));
 sky130_fd_sc_hd__mux4_2 _30620_ (.A0(_01110_),
    .A1(_01111_),
    .A2(_01112_),
    .A3(_01113_),
    .S0(net464),
    .S1(net472),
    .X(_01114_));
 sky130_fd_sc_hd__mux4_1 _30621_ (.A0(_01115_),
    .A1(_01116_),
    .A2(_01117_),
    .A3(_01118_),
    .S0(net464),
    .S1(net472),
    .X(_01119_));
 sky130_fd_sc_hd__mux4_2 _30622_ (.A0(_01104_),
    .A1(_01109_),
    .A2(_01114_),
    .A3(_01119_),
    .S0(net477),
    .S1(net480),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_1 _30623_ (.A0(_01094_),
    .A1(_01095_),
    .A2(_01096_),
    .A3(_01097_),
    .S0(net464),
    .S1(net472),
    .X(_01098_));
 sky130_fd_sc_hd__mux4_2 _30624_ (.A0(_01073_),
    .A1(_01074_),
    .A2(_01075_),
    .A3(_01076_),
    .S0(net464),
    .S1(net472),
    .X(_01077_));
 sky130_fd_sc_hd__mux4_2 _30625_ (.A0(_01078_),
    .A1(_01079_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(net464),
    .S1(net472),
    .X(_01082_));
 sky130_fd_sc_hd__mux4_2 _30626_ (.A0(_01083_),
    .A1(_01084_),
    .A2(_01085_),
    .A3(_01086_),
    .S0(net464),
    .S1(net472),
    .X(_01087_));
 sky130_fd_sc_hd__mux4_1 _30627_ (.A0(_01088_),
    .A1(_01089_),
    .A2(_01090_),
    .A3(_01091_),
    .S0(net464),
    .S1(net472),
    .X(_01092_));
 sky130_fd_sc_hd__mux4_1 _30628_ (.A0(_01077_),
    .A1(_01082_),
    .A2(_01087_),
    .A3(_01092_),
    .S0(net477),
    .S1(net480),
    .X(_01093_));
 sky130_fd_sc_hd__mux4_1 _30629_ (.A0(_01067_),
    .A1(_01068_),
    .A2(_01069_),
    .A3(_01070_),
    .S0(net465),
    .S1(net472),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_1 _30630_ (.A0(_01046_),
    .A1(_01047_),
    .A2(_01048_),
    .A3(_01049_),
    .S0(net465),
    .S1(net473),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_2 _30631_ (.A0(_01051_),
    .A1(_01052_),
    .A2(_01053_),
    .A3(_01054_),
    .S0(net465),
    .S1(net473),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_2 _30632_ (.A0(_01056_),
    .A1(_01057_),
    .A2(_01058_),
    .A3(_01059_),
    .S0(net465),
    .S1(net473),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_1 _30633_ (.A0(_01061_),
    .A1(_01062_),
    .A2(_01063_),
    .A3(_01064_),
    .S0(net465),
    .S1(net473),
    .X(_01065_));
 sky130_fd_sc_hd__mux4_2 _30634_ (.A0(_01050_),
    .A1(_01055_),
    .A2(_01060_),
    .A3(_01065_),
    .S0(net477),
    .S1(net480),
    .X(_01066_));
 sky130_fd_sc_hd__mux4_1 _30635_ (.A0(_01040_),
    .A1(_01041_),
    .A2(_01042_),
    .A3(_01043_),
    .S0(net467),
    .S1(net475),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_2 _30636_ (.A0(_01019_),
    .A1(_01020_),
    .A2(_01021_),
    .A3(_01022_),
    .S0(net467),
    .S1(net475),
    .X(_01023_));
 sky130_fd_sc_hd__mux4_2 _30637_ (.A0(_01024_),
    .A1(_01025_),
    .A2(_01026_),
    .A3(_01027_),
    .S0(net467),
    .S1(net475),
    .X(_01028_));
 sky130_fd_sc_hd__mux4_1 _30638_ (.A0(_01029_),
    .A1(_01030_),
    .A2(_01031_),
    .A3(_01032_),
    .S0(net467),
    .S1(net475),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_1 _30639_ (.A0(_01034_),
    .A1(_01035_),
    .A2(_01036_),
    .A3(_01037_),
    .S0(net467),
    .S1(net475),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_2 _30640_ (.A0(_01023_),
    .A1(_01028_),
    .A2(_01033_),
    .A3(_01038_),
    .S0(net477),
    .S1(net480),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_1 _30641_ (.A0(_01013_),
    .A1(_01014_),
    .A2(_01015_),
    .A3(_01016_),
    .S0(net465),
    .S1(net473),
    .X(_01017_));
 sky130_fd_sc_hd__mux4_1 _30642_ (.A0(_00992_),
    .A1(_00993_),
    .A2(_00994_),
    .A3(_00995_),
    .S0(net466),
    .S1(net473),
    .X(_00996_));
 sky130_fd_sc_hd__mux4_2 _30643_ (.A0(_00997_),
    .A1(_00998_),
    .A2(_00999_),
    .A3(_01000_),
    .S0(net466),
    .S1(net473),
    .X(_01001_));
 sky130_fd_sc_hd__mux4_2 _30644_ (.A0(_01002_),
    .A1(_01003_),
    .A2(_01004_),
    .A3(_01005_),
    .S0(net466),
    .S1(net473),
    .X(_01006_));
 sky130_fd_sc_hd__mux4_1 _30645_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(net466),
    .S1(net473),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_2 _30646_ (.A0(_00996_),
    .A1(_01001_),
    .A2(_01006_),
    .A3(_01011_),
    .S0(net477),
    .S1(net480),
    .X(_01012_));
 sky130_fd_sc_hd__mux4_1 _30647_ (.A0(_00986_),
    .A1(_00987_),
    .A2(_00988_),
    .A3(_00989_),
    .S0(net467),
    .S1(net475),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_2 _30648_ (.A0(_00965_),
    .A1(_00966_),
    .A2(_00967_),
    .A3(_00968_),
    .S0(net466),
    .S1(net475),
    .X(_00969_));
 sky130_fd_sc_hd__mux4_2 _30649_ (.A0(_00970_),
    .A1(_00971_),
    .A2(_00972_),
    .A3(_00973_),
    .S0(net467),
    .S1(net475),
    .X(_00974_));
 sky130_fd_sc_hd__mux4_1 _30650_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(net467),
    .S1(net475),
    .X(_00979_));
 sky130_fd_sc_hd__mux4_1 _30651_ (.A0(_00980_),
    .A1(_00981_),
    .A2(_00982_),
    .A3(_00983_),
    .S0(net466),
    .S1(net475),
    .X(_00984_));
 sky130_fd_sc_hd__mux4_2 _30652_ (.A0(_00969_),
    .A1(_00974_),
    .A2(_00979_),
    .A3(_00984_),
    .S0(net477),
    .S1(net480),
    .X(_00985_));
 sky130_fd_sc_hd__mux4_1 _30653_ (.A0(_00959_),
    .A1(_00960_),
    .A2(_00961_),
    .A3(_00962_),
    .S0(net465),
    .S1(net475),
    .X(_00963_));
 sky130_fd_sc_hd__mux4_2 _30654_ (.A0(_00938_),
    .A1(_00939_),
    .A2(_00940_),
    .A3(_00941_),
    .S0(net466),
    .S1(net473),
    .X(_00942_));
 sky130_fd_sc_hd__mux4_2 _30655_ (.A0(_00943_),
    .A1(_00944_),
    .A2(_00945_),
    .A3(_00946_),
    .S0(net466),
    .S1(net473),
    .X(_00947_));
 sky130_fd_sc_hd__mux4_1 _30656_ (.A0(_00948_),
    .A1(_00949_),
    .A2(_00950_),
    .A3(_00951_),
    .S0(net466),
    .S1(net473),
    .X(_00952_));
 sky130_fd_sc_hd__mux4_1 _30657_ (.A0(_00953_),
    .A1(_00954_),
    .A2(_00955_),
    .A3(_00956_),
    .S0(net466),
    .S1(net473),
    .X(_00957_));
 sky130_fd_sc_hd__mux4_2 _30658_ (.A0(_00942_),
    .A1(_00947_),
    .A2(_00952_),
    .A3(_00957_),
    .S0(net477),
    .S1(net480),
    .X(_00958_));
 sky130_fd_sc_hd__mux4_1 _30659_ (.A0(_00932_),
    .A1(_00933_),
    .A2(_00934_),
    .A3(_00935_),
    .S0(net466),
    .S1(net473),
    .X(_00936_));
 sky130_fd_sc_hd__mux4_2 _30660_ (.A0(_00911_),
    .A1(_00912_),
    .A2(_00913_),
    .A3(_00914_),
    .S0(net466),
    .S1(net473),
    .X(_00915_));
 sky130_fd_sc_hd__mux4_2 _30661_ (.A0(_00916_),
    .A1(_00917_),
    .A2(_00918_),
    .A3(_00919_),
    .S0(net466),
    .S1(net473),
    .X(_00920_));
 sky130_fd_sc_hd__mux4_1 _30662_ (.A0(_00921_),
    .A1(_00922_),
    .A2(_00923_),
    .A3(_00924_),
    .S0(net466),
    .S1(net473),
    .X(_00925_));
 sky130_fd_sc_hd__mux4_1 _30663_ (.A0(_00926_),
    .A1(_00927_),
    .A2(_00928_),
    .A3(_00929_),
    .S0(net466),
    .S1(net473),
    .X(_00930_));
 sky130_fd_sc_hd__mux4_2 _30664_ (.A0(_00915_),
    .A1(_00920_),
    .A2(_00925_),
    .A3(_00930_),
    .S0(net477),
    .S1(net480),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_1 _30665_ (.A0(_00905_),
    .A1(_00906_),
    .A2(_00907_),
    .A3(_00908_),
    .S0(net467),
    .S1(net475),
    .X(_00909_));
 sky130_fd_sc_hd__mux4_2 _30666_ (.A0(_00884_),
    .A1(_00885_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(net467),
    .S1(net475),
    .X(_00888_));
 sky130_fd_sc_hd__mux4_2 _30667_ (.A0(_00889_),
    .A1(_00890_),
    .A2(_00891_),
    .A3(_00892_),
    .S0(net467),
    .S1(net475),
    .X(_00893_));
 sky130_fd_sc_hd__mux4_1 _30668_ (.A0(_00894_),
    .A1(_00895_),
    .A2(_00896_),
    .A3(_00897_),
    .S0(net467),
    .S1(net475),
    .X(_00898_));
 sky130_fd_sc_hd__mux4_1 _30669_ (.A0(_00899_),
    .A1(_00900_),
    .A2(_00901_),
    .A3(_00902_),
    .S0(net467),
    .S1(net475),
    .X(_00903_));
 sky130_fd_sc_hd__mux4_2 _30670_ (.A0(_00888_),
    .A1(_00893_),
    .A2(_00898_),
    .A3(_00903_),
    .S0(net477),
    .S1(net480),
    .X(_00904_));
 sky130_fd_sc_hd__mux4_1 _30671_ (.A0(_00878_),
    .A1(_00879_),
    .A2(_00880_),
    .A3(_00881_),
    .S0(net459),
    .S1(net470),
    .X(_00882_));
 sky130_fd_sc_hd__mux4_2 _30672_ (.A0(_00857_),
    .A1(_00858_),
    .A2(_00859_),
    .A3(_00860_),
    .S0(net459),
    .S1(net470),
    .X(_00861_));
 sky130_fd_sc_hd__mux4_2 _30673_ (.A0(_00862_),
    .A1(_00863_),
    .A2(_00864_),
    .A3(_00865_),
    .S0(net459),
    .S1(net470),
    .X(_00866_));
 sky130_fd_sc_hd__mux4_2 _30674_ (.A0(_00867_),
    .A1(_00868_),
    .A2(_00869_),
    .A3(_00870_),
    .S0(net459),
    .S1(net470),
    .X(_00871_));
 sky130_fd_sc_hd__mux4_1 _30675_ (.A0(_00872_),
    .A1(_00873_),
    .A2(_00874_),
    .A3(_00875_),
    .S0(net459),
    .S1(net470),
    .X(_00876_));
 sky130_fd_sc_hd__mux4_2 _30676_ (.A0(_00861_),
    .A1(_00866_),
    .A2(_00871_),
    .A3(_00876_),
    .S0(net476),
    .S1(net479),
    .X(_00877_));
 sky130_fd_sc_hd__mux4_1 _30677_ (.A0(_00851_),
    .A1(_00852_),
    .A2(_00853_),
    .A3(_00854_),
    .S0(net461),
    .S1(net471),
    .X(_00855_));
 sky130_fd_sc_hd__mux4_2 _30678_ (.A0(_00830_),
    .A1(_00831_),
    .A2(_00832_),
    .A3(_00833_),
    .S0(net461),
    .S1(net471),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_2 _30679_ (.A0(_00835_),
    .A1(_00836_),
    .A2(_00837_),
    .A3(_00838_),
    .S0(net459),
    .S1(net470),
    .X(_00839_));
 sky130_fd_sc_hd__mux4_2 _30680_ (.A0(_00840_),
    .A1(_00841_),
    .A2(_00842_),
    .A3(_00843_),
    .S0(net461),
    .S1(net471),
    .X(_00844_));
 sky130_fd_sc_hd__mux4_1 _30681_ (.A0(_00845_),
    .A1(_00846_),
    .A2(_00847_),
    .A3(_00848_),
    .S0(net461),
    .S1(net471),
    .X(_00849_));
 sky130_fd_sc_hd__mux4_2 _30682_ (.A0(_00834_),
    .A1(_00839_),
    .A2(_00844_),
    .A3(_00849_),
    .S0(net478),
    .S1(net479),
    .X(_00850_));
 sky130_fd_sc_hd__mux4_1 _30683_ (.A0(_00824_),
    .A1(_00825_),
    .A2(_00826_),
    .A3(_00827_),
    .S0(net458),
    .S1(net469),
    .X(_00828_));
 sky130_fd_sc_hd__mux4_2 _30684_ (.A0(_00803_),
    .A1(_00804_),
    .A2(_00805_),
    .A3(_00806_),
    .S0(net461),
    .S1(net471),
    .X(_00807_));
 sky130_fd_sc_hd__mux4_2 _30685_ (.A0(_00808_),
    .A1(_00809_),
    .A2(_00810_),
    .A3(_00811_),
    .S0(net459),
    .S1(net469),
    .X(_00812_));
 sky130_fd_sc_hd__mux4_1 _30686_ (.A0(_00813_),
    .A1(_00814_),
    .A2(_00815_),
    .A3(_00816_),
    .S0(net461),
    .S1(net470),
    .X(_00817_));
 sky130_fd_sc_hd__mux4_1 _30687_ (.A0(_00818_),
    .A1(_00819_),
    .A2(_00820_),
    .A3(_00821_),
    .S0(net461),
    .S1(net471),
    .X(_00822_));
 sky130_fd_sc_hd__mux4_2 _30688_ (.A0(_00807_),
    .A1(_00812_),
    .A2(_00817_),
    .A3(_00822_),
    .S0(net476),
    .S1(net479),
    .X(_00823_));
 sky130_fd_sc_hd__mux4_1 _30689_ (.A0(_00797_),
    .A1(_00798_),
    .A2(_00799_),
    .A3(_00800_),
    .S0(net458),
    .S1(net469),
    .X(_00801_));
 sky130_fd_sc_hd__mux4_2 _30690_ (.A0(_00776_),
    .A1(_00777_),
    .A2(_00778_),
    .A3(_00779_),
    .S0(net461),
    .S1(net470),
    .X(_00780_));
 sky130_fd_sc_hd__mux4_2 _30691_ (.A0(_00781_),
    .A1(_00782_),
    .A2(_00783_),
    .A3(_00784_),
    .S0(net459),
    .S1(net469),
    .X(_00785_));
 sky130_fd_sc_hd__mux4_2 _30692_ (.A0(_00786_),
    .A1(_00787_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(net460),
    .S1(net470),
    .X(_00790_));
 sky130_fd_sc_hd__mux4_1 _30693_ (.A0(_00791_),
    .A1(_00792_),
    .A2(_00793_),
    .A3(_00794_),
    .S0(net461),
    .S1(net470),
    .X(_00795_));
 sky130_fd_sc_hd__mux4_2 _30694_ (.A0(_00780_),
    .A1(_00785_),
    .A2(_00790_),
    .A3(_00795_),
    .S0(net476),
    .S1(net479),
    .X(_00796_));
 sky130_fd_sc_hd__mux4_1 _30695_ (.A0(_00770_),
    .A1(_00771_),
    .A2(_00772_),
    .A3(_00773_),
    .S0(net460),
    .S1(net469),
    .X(_00774_));
 sky130_fd_sc_hd__mux4_1 _30696_ (.A0(_00749_),
    .A1(_00750_),
    .A2(_00751_),
    .A3(_00752_),
    .S0(net460),
    .S1(net469),
    .X(_00753_));
 sky130_fd_sc_hd__mux4_2 _30697_ (.A0(_00754_),
    .A1(_00755_),
    .A2(_00756_),
    .A3(_00757_),
    .S0(net459),
    .S1(net469),
    .X(_00758_));
 sky130_fd_sc_hd__mux4_2 _30698_ (.A0(_00759_),
    .A1(_00760_),
    .A2(_00761_),
    .A3(_00762_),
    .S0(net459),
    .S1(net470),
    .X(_00763_));
 sky130_fd_sc_hd__mux4_1 _30699_ (.A0(_00764_),
    .A1(_00765_),
    .A2(_00766_),
    .A3(_00767_),
    .S0(net459),
    .S1(net469),
    .X(_00768_));
 sky130_fd_sc_hd__mux4_2 _30700_ (.A0(_00753_),
    .A1(_00758_),
    .A2(_00763_),
    .A3(_00768_),
    .S0(net476),
    .S1(net479),
    .X(_00769_));
 sky130_fd_sc_hd__mux4_1 _30701_ (.A0(_00743_),
    .A1(_00744_),
    .A2(_00745_),
    .A3(_00746_),
    .S0(net461),
    .S1(net470),
    .X(_00747_));
 sky130_fd_sc_hd__mux4_2 _30702_ (.A0(_00722_),
    .A1(_00723_),
    .A2(_00724_),
    .A3(_00725_),
    .S0(net461),
    .S1(net470),
    .X(_00726_));
 sky130_fd_sc_hd__mux4_2 _30703_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(net459),
    .S1(net470),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_2 _30704_ (.A0(_00732_),
    .A1(_00733_),
    .A2(_00734_),
    .A3(_00735_),
    .S0(net461),
    .S1(net470),
    .X(_00736_));
 sky130_fd_sc_hd__mux4_1 _30705_ (.A0(_00737_),
    .A1(_00738_),
    .A2(_00739_),
    .A3(_00740_),
    .S0(net461),
    .S1(net470),
    .X(_00741_));
 sky130_fd_sc_hd__mux4_2 _30706_ (.A0(_00726_),
    .A1(_00731_),
    .A2(_00736_),
    .A3(_00741_),
    .S0(net476),
    .S1(net479),
    .X(_00742_));
 sky130_fd_sc_hd__mux4_2 _30707_ (.A0(_00716_),
    .A1(_00717_),
    .A2(_00718_),
    .A3(_00719_),
    .S0(net458),
    .S1(net469),
    .X(_00720_));
 sky130_fd_sc_hd__mux4_2 _30708_ (.A0(_00695_),
    .A1(_00696_),
    .A2(_00697_),
    .A3(_00698_),
    .S0(net458),
    .S1(net469),
    .X(_00699_));
 sky130_fd_sc_hd__mux4_2 _30709_ (.A0(_00700_),
    .A1(_00701_),
    .A2(_00702_),
    .A3(_00703_),
    .S0(net460),
    .S1(net469),
    .X(_00704_));
 sky130_fd_sc_hd__mux4_2 _30710_ (.A0(_00705_),
    .A1(_00706_),
    .A2(_00707_),
    .A3(_00708_),
    .S0(net458),
    .S1(net469),
    .X(_00709_));
 sky130_fd_sc_hd__mux4_1 _30711_ (.A0(_00710_),
    .A1(_00711_),
    .A2(_00712_),
    .A3(_00713_),
    .S0(net458),
    .S1(net469),
    .X(_00714_));
 sky130_fd_sc_hd__mux4_1 _30712_ (.A0(_00699_),
    .A1(_00704_),
    .A2(_00709_),
    .A3(_00714_),
    .S0(net476),
    .S1(net479),
    .X(_00715_));
 sky130_fd_sc_hd__mux4_1 _30713_ (.A0(_00689_),
    .A1(_00690_),
    .A2(_00691_),
    .A3(_00692_),
    .S0(net457),
    .S1(net468),
    .X(_00693_));
 sky130_fd_sc_hd__mux4_2 _30714_ (.A0(_00668_),
    .A1(_00669_),
    .A2(_00670_),
    .A3(_00671_),
    .S0(net457),
    .S1(net468),
    .X(_00672_));
 sky130_fd_sc_hd__mux4_2 _30715_ (.A0(_00673_),
    .A1(_00674_),
    .A2(_00675_),
    .A3(_00676_),
    .S0(net457),
    .S1(net468),
    .X(_00677_));
 sky130_fd_sc_hd__mux4_1 _30716_ (.A0(_00678_),
    .A1(_00679_),
    .A2(_00680_),
    .A3(_00681_),
    .S0(net457),
    .S1(net468),
    .X(_00682_));
 sky130_fd_sc_hd__mux4_1 _30717_ (.A0(_00683_),
    .A1(_00684_),
    .A2(_00685_),
    .A3(_00686_),
    .S0(net457),
    .S1(net468),
    .X(_00687_));
 sky130_fd_sc_hd__mux4_2 _30718_ (.A0(_00672_),
    .A1(_00677_),
    .A2(_00682_),
    .A3(_00687_),
    .S0(net476),
    .S1(net479),
    .X(_00688_));
 sky130_fd_sc_hd__mux4_1 _30719_ (.A0(_00662_),
    .A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .S0(net460),
    .S1(net468),
    .X(_00666_));
 sky130_fd_sc_hd__mux4_1 _30720_ (.A0(_00641_),
    .A1(_00642_),
    .A2(_00643_),
    .A3(_00644_),
    .S0(net457),
    .S1(net468),
    .X(_00645_));
 sky130_fd_sc_hd__mux4_2 _30721_ (.A0(_00646_),
    .A1(_00647_),
    .A2(_00648_),
    .A3(_00649_),
    .S0(net457),
    .S1(net468),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_1 _30722_ (.A0(_00651_),
    .A1(_00652_),
    .A2(_00653_),
    .A3(_00654_),
    .S0(net457),
    .S1(net468),
    .X(_00655_));
 sky130_fd_sc_hd__mux4_2 _30723_ (.A0(_00656_),
    .A1(_00657_),
    .A2(_00658_),
    .A3(_00659_),
    .S0(net457),
    .S1(net468),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_2 _30724_ (.A0(_00645_),
    .A1(_00650_),
    .A2(_00655_),
    .A3(_00660_),
    .S0(net476),
    .S1(net479),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_1 _30725_ (.A0(_00635_),
    .A1(_00636_),
    .A2(_00637_),
    .A3(_00638_),
    .S0(net457),
    .S1(net468),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_1 _30726_ (.A0(_00614_),
    .A1(_00615_),
    .A2(_00616_),
    .A3(_00617_),
    .S0(net460),
    .S1(net468),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_2 _30727_ (.A0(_00619_),
    .A1(_00620_),
    .A2(_00621_),
    .A3(_00622_),
    .S0(net457),
    .S1(net468),
    .X(_00623_));
 sky130_fd_sc_hd__mux4_1 _30728_ (.A0(_00624_),
    .A1(_00625_),
    .A2(_00626_),
    .A3(_00627_),
    .S0(net460),
    .S1(net468),
    .X(_00628_));
 sky130_fd_sc_hd__mux4_2 _30729_ (.A0(_00629_),
    .A1(_00630_),
    .A2(_00631_),
    .A3(_00632_),
    .S0(net457),
    .S1(net468),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_1 _30730_ (.A0(_00618_),
    .A1(_00623_),
    .A2(_00628_),
    .A3(_00633_),
    .S0(net476),
    .S1(net479),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_1 _30731_ (.A0(_00608_),
    .A1(_00609_),
    .A2(_00610_),
    .A3(_00611_),
    .S0(net460),
    .S1(net468),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_2 _30732_ (.A0(_00587_),
    .A1(_00588_),
    .A2(_00589_),
    .A3(_00590_),
    .S0(net458),
    .S1(net469),
    .X(_00591_));
 sky130_fd_sc_hd__mux4_2 _30733_ (.A0(_00592_),
    .A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .S0(net460),
    .S1(net468),
    .X(_00596_));
 sky130_fd_sc_hd__mux4_1 _30734_ (.A0(_00597_),
    .A1(_00598_),
    .A2(_00599_),
    .A3(_00600_),
    .S0(net458),
    .S1(net468),
    .X(_00601_));
 sky130_fd_sc_hd__mux4_2 _30735_ (.A0(_00602_),
    .A1(_00603_),
    .A2(_00604_),
    .A3(_00605_),
    .S0(net460),
    .S1(net468),
    .X(_00606_));
 sky130_fd_sc_hd__mux4_2 _30736_ (.A0(_00591_),
    .A1(_00596_),
    .A2(_00601_),
    .A3(_00606_),
    .S0(net476),
    .S1(net479),
    .X(_00607_));
 sky130_fd_sc_hd__mux4_1 _30737_ (.A0(_00581_),
    .A1(_00582_),
    .A2(_00583_),
    .A3(_00584_),
    .S0(net457),
    .S1(net468),
    .X(_00585_));
 sky130_fd_sc_hd__mux4_1 _30738_ (.A0(_00560_),
    .A1(_00561_),
    .A2(_00562_),
    .A3(_00563_),
    .S0(net457),
    .S1(net468),
    .X(_00564_));
 sky130_fd_sc_hd__mux4_2 _30739_ (.A0(_00565_),
    .A1(_00566_),
    .A2(_00567_),
    .A3(_00568_),
    .S0(net457),
    .S1(net468),
    .X(_00569_));
 sky130_fd_sc_hd__mux4_1 _30740_ (.A0(_00570_),
    .A1(_00571_),
    .A2(_00572_),
    .A3(_00573_),
    .S0(net457),
    .S1(net468),
    .X(_00574_));
 sky130_fd_sc_hd__mux4_2 _30741_ (.A0(_00575_),
    .A1(_00576_),
    .A2(_00577_),
    .A3(_00578_),
    .S0(net457),
    .S1(net468),
    .X(_00579_));
 sky130_fd_sc_hd__mux4_2 _30742_ (.A0(_00564_),
    .A1(_00569_),
    .A2(_00574_),
    .A3(_00579_),
    .S0(net476),
    .S1(net479),
    .X(_00580_));
 sky130_fd_sc_hd__mux4_1 _30743_ (.A0(_00554_),
    .A1(_00555_),
    .A2(_00556_),
    .A3(_00557_),
    .S0(net462),
    .S1(net471),
    .X(_00558_));
 sky130_fd_sc_hd__mux4_2 _30744_ (.A0(_00533_),
    .A1(_00534_),
    .A2(_00535_),
    .A3(_00536_),
    .S0(net462),
    .S1(net471),
    .X(_00537_));
 sky130_fd_sc_hd__mux4_2 _30745_ (.A0(_00538_),
    .A1(_00539_),
    .A2(_00540_),
    .A3(_00541_),
    .S0(net461),
    .S1(net471),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_1 _30746_ (.A0(_00543_),
    .A1(_00544_),
    .A2(_00545_),
    .A3(_00546_),
    .S0(net461),
    .S1(net471),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_2 _30747_ (.A0(_00548_),
    .A1(_00549_),
    .A2(_00550_),
    .A3(_00551_),
    .S0(net462),
    .S1(net471),
    .X(_00552_));
 sky130_fd_sc_hd__mux4_2 _30748_ (.A0(_00537_),
    .A1(_00542_),
    .A2(_00547_),
    .A3(_00552_),
    .S0(net478),
    .S1(net479),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_1 _30749_ (.A0(_00527_),
    .A1(_00528_),
    .A2(_00529_),
    .A3(_00530_),
    .S0(net462),
    .S1(net471),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_2 _30750_ (.A0(_00506_),
    .A1(_00507_),
    .A2(_00508_),
    .A3(_00509_),
    .S0(net462),
    .S1(net474),
    .X(_00510_));
 sky130_fd_sc_hd__mux4_2 _30751_ (.A0(_00511_),
    .A1(_00512_),
    .A2(_00513_),
    .A3(_00514_),
    .S0(net462),
    .S1(net471),
    .X(_00515_));
 sky130_fd_sc_hd__mux4_2 _30752_ (.A0(_00516_),
    .A1(_00517_),
    .A2(_00518_),
    .A3(_00519_),
    .S0(net462),
    .S1(net471),
    .X(_00520_));
 sky130_fd_sc_hd__mux4_1 _30753_ (.A0(_00521_),
    .A1(_00522_),
    .A2(_00523_),
    .A3(_00524_),
    .S0(net462),
    .S1(net471),
    .X(_00525_));
 sky130_fd_sc_hd__mux4_2 _30754_ (.A0(_00510_),
    .A1(_00515_),
    .A2(_00520_),
    .A3(_00525_),
    .S0(net478),
    .S1(net479),
    .X(_00526_));
 sky130_fd_sc_hd__mux4_1 _30755_ (.A0(_00500_),
    .A1(_00501_),
    .A2(_00502_),
    .A3(_00503_),
    .S0(net462),
    .S1(net471),
    .X(_00504_));
 sky130_fd_sc_hd__mux4_2 _30756_ (.A0(_00479_),
    .A1(_00480_),
    .A2(_00481_),
    .A3(_00482_),
    .S0(net462),
    .S1(net471),
    .X(_00483_));
 sky130_fd_sc_hd__mux4_2 _30757_ (.A0(_00484_),
    .A1(_00485_),
    .A2(_00486_),
    .A3(_00487_),
    .S0(net462),
    .S1(net471),
    .X(_00488_));
 sky130_fd_sc_hd__mux4_2 _30758_ (.A0(_00489_),
    .A1(_00490_),
    .A2(_00491_),
    .A3(_00492_),
    .S0(net462),
    .S1(net471),
    .X(_00493_));
 sky130_fd_sc_hd__mux4_1 _30759_ (.A0(_00494_),
    .A1(_00495_),
    .A2(_00496_),
    .A3(_00497_),
    .S0(net462),
    .S1(net471),
    .X(_00498_));
 sky130_fd_sc_hd__mux4_2 _30760_ (.A0(_00483_),
    .A1(_00488_),
    .A2(_00493_),
    .A3(_00498_),
    .S0(net478),
    .S1(net479),
    .X(_00499_));
 sky130_fd_sc_hd__mux4_1 _30761_ (.A0(_00473_),
    .A1(_00474_),
    .A2(_00475_),
    .A3(_00476_),
    .S0(net463),
    .S1(net474),
    .X(_00477_));
 sky130_fd_sc_hd__mux4_2 _30762_ (.A0(_00452_),
    .A1(_00453_),
    .A2(_00454_),
    .A3(_00455_),
    .S0(net463),
    .S1(net474),
    .X(_00456_));
 sky130_fd_sc_hd__mux4_2 _30763_ (.A0(_00457_),
    .A1(_00458_),
    .A2(_00459_),
    .A3(_00460_),
    .S0(net463),
    .S1(net474),
    .X(_00461_));
 sky130_fd_sc_hd__mux4_2 _30764_ (.A0(_00462_),
    .A1(_00463_),
    .A2(_00464_),
    .A3(_00465_),
    .S0(net463),
    .S1(net474),
    .X(_00466_));
 sky130_fd_sc_hd__mux4_1 _30765_ (.A0(_00467_),
    .A1(_00468_),
    .A2(_00469_),
    .A3(_00470_),
    .S0(net463),
    .S1(net474),
    .X(_00471_));
 sky130_fd_sc_hd__mux4_2 _30766_ (.A0(_00456_),
    .A1(_00461_),
    .A2(_00466_),
    .A3(_00471_),
    .S0(net478),
    .S1(_00362_),
    .X(_00472_));
 sky130_fd_sc_hd__mux4_1 _30767_ (.A0(_00446_),
    .A1(_00447_),
    .A2(_00448_),
    .A3(_00449_),
    .S0(net463),
    .S1(net474),
    .X(_00450_));
 sky130_fd_sc_hd__mux4_2 _30768_ (.A0(_00425_),
    .A1(_00426_),
    .A2(_00427_),
    .A3(_00428_),
    .S0(net463),
    .S1(net474),
    .X(_00429_));
 sky130_fd_sc_hd__mux4_2 _30769_ (.A0(_00430_),
    .A1(_00431_),
    .A2(_00432_),
    .A3(_00433_),
    .S0(net463),
    .S1(net474),
    .X(_00434_));
 sky130_fd_sc_hd__mux4_2 _30770_ (.A0(_00435_),
    .A1(_00436_),
    .A2(_00437_),
    .A3(_00438_),
    .S0(net463),
    .S1(net474),
    .X(_00439_));
 sky130_fd_sc_hd__mux4_1 _30771_ (.A0(_00440_),
    .A1(_00441_),
    .A2(_00442_),
    .A3(_00443_),
    .S0(net463),
    .S1(net474),
    .X(_00444_));
 sky130_fd_sc_hd__mux4_2 _30772_ (.A0(_00429_),
    .A1(_00434_),
    .A2(_00439_),
    .A3(_00444_),
    .S0(net478),
    .S1(_00362_),
    .X(_00445_));
 sky130_fd_sc_hd__mux4_2 _30773_ (.A0(_00419_),
    .A1(_00420_),
    .A2(_00421_),
    .A3(_00422_),
    .S0(net463),
    .S1(net474),
    .X(_00423_));
 sky130_fd_sc_hd__mux4_1 _30774_ (.A0(_00398_),
    .A1(_00399_),
    .A2(_00400_),
    .A3(_00401_),
    .S0(net463),
    .S1(net474),
    .X(_00402_));
 sky130_fd_sc_hd__mux4_2 _30775_ (.A0(_00403_),
    .A1(_00404_),
    .A2(_00405_),
    .A3(_00406_),
    .S0(net463),
    .S1(net474),
    .X(_00407_));
 sky130_fd_sc_hd__mux4_1 _30776_ (.A0(_00408_),
    .A1(_00409_),
    .A2(_00410_),
    .A3(_00411_),
    .S0(net463),
    .S1(net474),
    .X(_00412_));
 sky130_fd_sc_hd__mux4_2 _30777_ (.A0(_00413_),
    .A1(_00414_),
    .A2(_00415_),
    .A3(_00416_),
    .S0(net463),
    .S1(net474),
    .X(_00417_));
 sky130_fd_sc_hd__mux4_2 _30778_ (.A0(_00402_),
    .A1(_00407_),
    .A2(_00412_),
    .A3(_00417_),
    .S0(net478),
    .S1(_00362_),
    .X(_00418_));
 sky130_fd_sc_hd__mux4_1 _30779_ (.A0(_00392_),
    .A1(_00393_),
    .A2(_00394_),
    .A3(_00395_),
    .S0(net458),
    .S1(net469),
    .X(_00396_));
 sky130_fd_sc_hd__mux4_2 _30780_ (.A0(_00371_),
    .A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .S0(net462),
    .S1(net471),
    .X(_00375_));
 sky130_fd_sc_hd__mux4_1 _30781_ (.A0(_00376_),
    .A1(_00377_),
    .A2(_00378_),
    .A3(_00379_),
    .S0(net458),
    .S1(net469),
    .X(_00380_));
 sky130_fd_sc_hd__mux4_2 _30782_ (.A0(_00381_),
    .A1(_00382_),
    .A2(_00383_),
    .A3(_00384_),
    .S0(net458),
    .S1(net469),
    .X(_00385_));
 sky130_fd_sc_hd__mux4_1 _30783_ (.A0(_00386_),
    .A1(_00387_),
    .A2(_00388_),
    .A3(_00389_),
    .S0(net458),
    .S1(net469),
    .X(_00390_));
 sky130_fd_sc_hd__mux4_2 _30784_ (.A0(_00375_),
    .A1(_00380_),
    .A2(_00385_),
    .A3(_00390_),
    .S0(net476),
    .S1(net479),
    .X(_00391_));
 sky130_fd_sc_hd__mux4_1 _30785_ (.A0(\cpuregs[16][0] ),
    .A1(\cpuregs[17][0] ),
    .A2(\cpuregs[18][0] ),
    .A3(\cpuregs[19][0] ),
    .S0(_00357_),
    .S1(net475),
    .X(_00369_));
 sky130_fd_sc_hd__mux4_2 _30786_ (.A0(\cpuregs[0][0] ),
    .A1(\cpuregs[1][0] ),
    .A2(\cpuregs[2][0] ),
    .A3(\cpuregs[3][0] ),
    .S0(_00357_),
    .S1(net475),
    .X(_00359_));
 sky130_fd_sc_hd__mux4_2 _30787_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .A2(\cpuregs[6][0] ),
    .A3(\cpuregs[7][0] ),
    .S0(net467),
    .S1(net474),
    .X(_00361_));
 sky130_fd_sc_hd__mux4_1 _30788_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .A2(\cpuregs[10][0] ),
    .A3(\cpuregs[11][0] ),
    .S0(net467),
    .S1(net474),
    .X(_00363_));
 sky130_fd_sc_hd__mux4_1 _30789_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .A2(\cpuregs[14][0] ),
    .A3(\cpuregs[15][0] ),
    .S0(_00357_),
    .S1(net474),
    .X(_00364_));
 sky130_fd_sc_hd__mux4_2 _30790_ (.A0(_00359_),
    .A1(_00361_),
    .A2(_00363_),
    .A3(_00364_),
    .S0(net478),
    .S1(net480),
    .X(_00365_));
 sky130_fd_sc_hd__mux4_1 _30791_ (.A0(_02581_),
    .A1(_01681_),
    .A2(_01679_),
    .A3(_02581_),
    .S0(net426),
    .S1(_00309_),
    .X(_01682_));
 sky130_fd_sc_hd__mux4_1 _30792_ (.A0(_02580_),
    .A1(_01677_),
    .A2(_01675_),
    .A3(_02580_),
    .S0(net426),
    .S1(_00309_),
    .X(_01678_));
 sky130_fd_sc_hd__mux4_1 _30793_ (.A0(_02579_),
    .A1(_01673_),
    .A2(_01671_),
    .A3(_02579_),
    .S0(net426),
    .S1(_00309_),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_2 _30794_ (.A0(_02578_),
    .A1(_01669_),
    .A2(_01667_),
    .A3(_02578_),
    .S0(net426),
    .S1(_00309_),
    .X(_01670_));
 sky130_fd_sc_hd__mux4_1 _30795_ (.A0(_02577_),
    .A1(_01665_),
    .A2(_01663_),
    .A3(_02577_),
    .S0(net426),
    .S1(_00309_),
    .X(_01666_));
 sky130_fd_sc_hd__mux4_1 _30796_ (.A0(_02576_),
    .A1(_01661_),
    .A2(_01659_),
    .A3(_02576_),
    .S0(net426),
    .S1(_00309_),
    .X(_01662_));
 sky130_fd_sc_hd__mux4_1 _30797_ (.A0(_02575_),
    .A1(_01657_),
    .A2(_01655_),
    .A3(_02575_),
    .S0(net426),
    .S1(_00309_),
    .X(_01658_));
 sky130_fd_sc_hd__mux4_1 _30798_ (.A0(_02574_),
    .A1(_01653_),
    .A2(_01651_),
    .A3(_02574_),
    .S0(net426),
    .S1(_00309_),
    .X(_01654_));
 sky130_fd_sc_hd__mux4_2 _30799_ (.A0(_02573_),
    .A1(_01649_),
    .A2(_01647_),
    .A3(_02573_),
    .S0(net426),
    .S1(_00309_),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_2 _30800_ (.A0(_02572_),
    .A1(_01645_),
    .A2(_01643_),
    .A3(_02572_),
    .S0(net426),
    .S1(_00309_),
    .X(_01646_));
 sky130_fd_sc_hd__mux4_1 _30801_ (.A0(_02570_),
    .A1(_01641_),
    .A2(_01639_),
    .A3(_02570_),
    .S0(net426),
    .S1(_00309_),
    .X(_01642_));
 sky130_fd_sc_hd__mux4_1 _30802_ (.A0(_02569_),
    .A1(_01637_),
    .A2(_01635_),
    .A3(_02569_),
    .S0(net426),
    .S1(_00309_),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_1 _30803_ (.A0(_02568_),
    .A1(_01633_),
    .A2(_01631_),
    .A3(_02568_),
    .S0(net426),
    .S1(_00309_),
    .X(_01634_));
 sky130_fd_sc_hd__mux4_1 _30804_ (.A0(_02567_),
    .A1(_01629_),
    .A2(_01627_),
    .A3(_02567_),
    .S0(net426),
    .S1(_00309_),
    .X(_01630_));
 sky130_fd_sc_hd__mux4_1 _30805_ (.A0(_02566_),
    .A1(_01625_),
    .A2(_01623_),
    .A3(_02566_),
    .S0(net426),
    .S1(_00309_),
    .X(_01626_));
 sky130_fd_sc_hd__mux4_1 _30806_ (.A0(_02565_),
    .A1(_01621_),
    .A2(_01619_),
    .A3(_02565_),
    .S0(net426),
    .S1(_00309_),
    .X(_01622_));
 sky130_fd_sc_hd__mux4_1 _30807_ (.A0(_02564_),
    .A1(_01617_),
    .A2(_01615_),
    .A3(_02564_),
    .S0(net426),
    .S1(_00309_),
    .X(_01618_));
 sky130_fd_sc_hd__mux4_1 _30808_ (.A0(_02563_),
    .A1(_01613_),
    .A2(_01611_),
    .A3(_02563_),
    .S0(net426),
    .S1(_00309_),
    .X(_01614_));
 sky130_fd_sc_hd__mux4_1 _30809_ (.A0(_02562_),
    .A1(_01609_),
    .A2(_01607_),
    .A3(_02562_),
    .S0(net426),
    .S1(_00309_),
    .X(_01610_));
 sky130_fd_sc_hd__mux4_1 _30810_ (.A0(_02561_),
    .A1(_01605_),
    .A2(_01603_),
    .A3(_02561_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01606_));
 sky130_fd_sc_hd__mux4_1 _30811_ (.A0(_02589_),
    .A1(_01601_),
    .A2(_01599_),
    .A3(_02589_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01602_));
 sky130_fd_sc_hd__mux4_1 _30812_ (.A0(_02588_),
    .A1(_01597_),
    .A2(_01595_),
    .A3(_02588_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01598_));
 sky130_fd_sc_hd__mux4_1 _30813_ (.A0(_02587_),
    .A1(_01593_),
    .A2(_01591_),
    .A3(_02587_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01594_));
 sky130_fd_sc_hd__mux4_1 _30814_ (.A0(_02586_),
    .A1(_01589_),
    .A2(_01587_),
    .A3(_02586_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _30815_ (.A0(_02585_),
    .A1(_01585_),
    .A2(_01583_),
    .A3(_02585_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01586_));
 sky130_fd_sc_hd__mux4_1 _30816_ (.A0(_02584_),
    .A1(_01581_),
    .A2(_01579_),
    .A3(_02584_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01582_));
 sky130_fd_sc_hd__mux4_1 _30817_ (.A0(_02583_),
    .A1(_01577_),
    .A2(_01575_),
    .A3(_02583_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01578_));
 sky130_fd_sc_hd__mux4_1 _30818_ (.A0(_02582_),
    .A1(_01573_),
    .A2(_01571_),
    .A3(_02582_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01574_));
 sky130_fd_sc_hd__mux4_1 _30819_ (.A0(_02571_),
    .A1(_01569_),
    .A2(_01567_),
    .A3(_02571_),
    .S0(_15209_),
    .S1(_00309_),
    .X(_01570_));
 sky130_fd_sc_hd__dfxtp_1 _30820_ (.D(_02687_),
    .Q(\alu_shl[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30821_ (.D(_02688_),
    .Q(\alu_shl[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30822_ (.D(_02689_),
    .Q(\alu_shl[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30823_ (.D(_02690_),
    .Q(\alu_shl[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30824_ (.D(_02691_),
    .Q(\alu_shl[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30825_ (.D(_02692_),
    .Q(\alu_shl[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30826_ (.D(_02693_),
    .Q(\alu_shl[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30827_ (.D(_02694_),
    .Q(\alu_shl[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30828_ (.D(_02695_),
    .Q(\alu_shl[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30829_ (.D(_02696_),
    .Q(\alu_shl[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30830_ (.D(_02697_),
    .Q(\alu_shl[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30831_ (.D(_02698_),
    .Q(\alu_shl[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30832_ (.D(_02699_),
    .Q(\alu_shl[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30833_ (.D(_02700_),
    .Q(\alu_shl[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30834_ (.D(_02701_),
    .Q(\alu_shl[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30835_ (.D(_02702_),
    .Q(\alu_shl[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30836_ (.D(_02703_),
    .Q(alu_wait),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30837_ (.D(_02704_),
    .Q(\latched_rd[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30838_ (.D(_02705_),
    .Q(\latched_rd[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30839_ (.D(_02706_),
    .Q(\latched_rd[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30840_ (.D(_02707_),
    .Q(\latched_rd[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30841_ (.D(_02708_),
    .Q(\decoded_imm[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30842_ (.D(_02709_),
    .Q(\decoded_imm[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30843_ (.D(_02710_),
    .Q(\decoded_imm[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30844_ (.D(_02711_),
    .Q(\decoded_imm[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30845_ (.D(_02712_),
    .Q(\decoded_imm[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30846_ (.D(_02713_),
    .Q(\decoded_imm[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30847_ (.D(_02714_),
    .Q(\decoded_imm[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30848_ (.D(_02715_),
    .Q(\decoded_imm[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30849_ (.D(_02716_),
    .Q(\decoded_imm[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30850_ (.D(_02717_),
    .Q(\decoded_imm[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30851_ (.D(_02718_),
    .Q(\decoded_imm[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30852_ (.D(_02719_),
    .Q(\decoded_imm[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30853_ (.D(_02720_),
    .Q(\decoded_imm[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30854_ (.D(_02721_),
    .Q(\decoded_imm[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30855_ (.D(_02722_),
    .Q(\decoded_imm[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30856_ (.D(_02723_),
    .Q(\decoded_imm[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30857_ (.D(_02724_),
    .Q(\decoded_imm[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30858_ (.D(_02725_),
    .Q(\decoded_imm[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30859_ (.D(_02726_),
    .Q(\decoded_imm[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30860_ (.D(_02727_),
    .Q(\decoded_imm[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30861_ (.D(_02728_),
    .Q(\decoded_imm[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30862_ (.D(_02729_),
    .Q(\decoded_imm[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30863_ (.D(_02730_),
    .Q(\decoded_imm[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30864_ (.D(_02731_),
    .Q(\decoded_imm[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30865_ (.D(_02732_),
    .Q(\decoded_imm[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30866_ (.D(_02733_),
    .Q(\decoded_imm[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30867_ (.D(_02734_),
    .Q(\decoded_imm[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30868_ (.D(_02735_),
    .Q(\decoded_imm[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30869_ (.D(_02736_),
    .Q(\decoded_imm[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30870_ (.D(_02737_),
    .Q(\decoded_imm[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30871_ (.D(_02738_),
    .Q(\decoded_imm[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30872_ (.D(_02739_),
    .Q(\irq_pending[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30873_ (.D(_02740_),
    .Q(\irq_pending[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30874_ (.D(_02741_),
    .Q(\irq_pending[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30875_ (.D(_02742_),
    .Q(\irq_pending[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30876_ (.D(_02743_),
    .Q(\irq_pending[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30877_ (.D(_02744_),
    .Q(\irq_pending[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30878_ (.D(_02745_),
    .Q(\irq_pending[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30879_ (.D(_02746_),
    .Q(\irq_pending[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30880_ (.D(_02747_),
    .Q(\irq_pending[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30881_ (.D(_02748_),
    .Q(\irq_pending[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30882_ (.D(_02749_),
    .Q(\irq_pending[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30883_ (.D(_02750_),
    .Q(\irq_pending[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30884_ (.D(_02751_),
    .Q(\irq_pending[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30885_ (.D(_02752_),
    .Q(\irq_pending[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30886_ (.D(_02753_),
    .Q(\irq_pending[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30887_ (.D(_02754_),
    .Q(\irq_pending[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30888_ (.D(_02755_),
    .Q(\irq_pending[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30889_ (.D(_02756_),
    .Q(\irq_pending[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30890_ (.D(_02757_),
    .Q(\irq_pending[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30891_ (.D(_02758_),
    .Q(\irq_pending[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30892_ (.D(_02759_),
    .Q(\irq_pending[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30893_ (.D(_02760_),
    .Q(\irq_pending[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30894_ (.D(_02761_),
    .Q(\irq_pending[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30895_ (.D(_02762_),
    .Q(\irq_pending[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30896_ (.D(_02763_),
    .Q(\irq_pending[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30897_ (.D(_02764_),
    .Q(\irq_pending[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30898_ (.D(_02765_),
    .Q(\irq_pending[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30899_ (.D(_02766_),
    .Q(\irq_pending[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30900_ (.D(_02767_),
    .Q(\irq_pending[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30901_ (.D(_02768_),
    .Q(\irq_pending[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30902_ (.D(_02769_),
    .Q(\irq_pending[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30903_ (.D(_02770_),
    .Q(\reg_next_pc[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30904_ (.D(_00045_),
    .Q(\mem_wordsize[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30905_ (.D(_00046_),
    .Q(\mem_wordsize[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30906_ (.D(_00047_),
    .Q(\mem_wordsize[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30907_ (.D(_15211_),
    .Q(\reg_out[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30908_ (.D(_15222_),
    .Q(\reg_out[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30909_ (.D(_15233_),
    .Q(\reg_out[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30910_ (.D(_15236_),
    .Q(\reg_out[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30911_ (.D(_15237_),
    .Q(\reg_out[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30912_ (.D(_15238_),
    .Q(\reg_out[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30913_ (.D(_15239_),
    .Q(\reg_out[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30914_ (.D(_15240_),
    .Q(\reg_out[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30915_ (.D(_15241_),
    .Q(\reg_out[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30916_ (.D(_15242_),
    .Q(\reg_out[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30917_ (.D(_15212_),
    .Q(\reg_out[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30918_ (.D(_15213_),
    .Q(\reg_out[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30919_ (.D(_15214_),
    .Q(\reg_out[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30920_ (.D(_15215_),
    .Q(\reg_out[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30921_ (.D(_15216_),
    .Q(\reg_out[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30922_ (.D(_15217_),
    .Q(\reg_out[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30923_ (.D(_15218_),
    .Q(\reg_out[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30924_ (.D(_15219_),
    .Q(\reg_out[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30925_ (.D(_15220_),
    .Q(\reg_out[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30926_ (.D(_15221_),
    .Q(\reg_out[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30927_ (.D(_15223_),
    .Q(\reg_out[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30928_ (.D(_15224_),
    .Q(\reg_out[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30929_ (.D(_15225_),
    .Q(\reg_out[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30930_ (.D(_15226_),
    .Q(\reg_out[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30931_ (.D(_15227_),
    .Q(\reg_out[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30932_ (.D(_15228_),
    .Q(\reg_out[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30933_ (.D(_15229_),
    .Q(\reg_out[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30934_ (.D(_15230_),
    .Q(\reg_out[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30935_ (.D(_15231_),
    .Q(\reg_out[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30936_ (.D(_15232_),
    .Q(\reg_out[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30937_ (.D(_15234_),
    .Q(\reg_out[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30938_ (.D(_15235_),
    .Q(\reg_out[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30939_ (.D(_00004_),
    .Q(\irq_pending[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30940_ (.D(_00003_),
    .Q(decoder_trigger),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30941_ (.D(\alu_out[0] ),
    .Q(\alu_out_q[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30942_ (.D(\alu_out[1] ),
    .Q(\alu_out_q[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30943_ (.D(\alu_out[2] ),
    .Q(\alu_out_q[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30944_ (.D(\alu_out[3] ),
    .Q(\alu_out_q[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30945_ (.D(\alu_out[4] ),
    .Q(\alu_out_q[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30946_ (.D(\alu_out[5] ),
    .Q(\alu_out_q[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30947_ (.D(\alu_out[6] ),
    .Q(\alu_out_q[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30948_ (.D(\alu_out[7] ),
    .Q(\alu_out_q[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30949_ (.D(\alu_out[8] ),
    .Q(\alu_out_q[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30950_ (.D(\alu_out[9] ),
    .Q(\alu_out_q[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30951_ (.D(\alu_out[10] ),
    .Q(\alu_out_q[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30952_ (.D(\alu_out[11] ),
    .Q(\alu_out_q[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30953_ (.D(\alu_out[12] ),
    .Q(\alu_out_q[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30954_ (.D(\alu_out[13] ),
    .Q(\alu_out_q[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30955_ (.D(\alu_out[14] ),
    .Q(\alu_out_q[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30956_ (.D(\alu_out[15] ),
    .Q(\alu_out_q[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30957_ (.D(\alu_out[16] ),
    .Q(\alu_out_q[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30958_ (.D(\alu_out[17] ),
    .Q(\alu_out_q[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30959_ (.D(\alu_out[18] ),
    .Q(\alu_out_q[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30960_ (.D(\alu_out[19] ),
    .Q(\alu_out_q[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30961_ (.D(\alu_out[20] ),
    .Q(\alu_out_q[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30962_ (.D(\alu_out[21] ),
    .Q(\alu_out_q[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30963_ (.D(\alu_out[22] ),
    .Q(\alu_out_q[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30964_ (.D(\alu_out[23] ),
    .Q(\alu_out_q[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30965_ (.D(\alu_out[24] ),
    .Q(\alu_out_q[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30966_ (.D(\alu_out[25] ),
    .Q(\alu_out_q[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30967_ (.D(\alu_out[26] ),
    .Q(\alu_out_q[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30968_ (.D(\alu_out[27] ),
    .Q(\alu_out_q[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30969_ (.D(\alu_out[28] ),
    .Q(\alu_out_q[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30970_ (.D(\alu_out[29] ),
    .Q(\alu_out_q[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30971_ (.D(\alu_out[30] ),
    .Q(\alu_out_q[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _30972_ (.D(\alu_out[31] ),
    .Q(\alu_out_q[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _30973_ (.D(_00005_),
    .Q(is_lui_auipc_jal),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30974_ (.D(_00006_),
    .Q(is_slti_blt_slt),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30975_ (.D(_00007_),
    .Q(is_sltiu_bltu_sltu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30976_ (.D(_02591_),
    .Q(\alu_add_sub[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30977_ (.D(_02602_),
    .Q(\alu_add_sub[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30978_ (.D(_02613_),
    .Q(\alu_add_sub[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30979_ (.D(_02616_),
    .Q(\alu_add_sub[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30980_ (.D(_02617_),
    .Q(\alu_add_sub[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30981_ (.D(_02618_),
    .Q(\alu_add_sub[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30982_ (.D(_02619_),
    .Q(\alu_add_sub[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30983_ (.D(_02620_),
    .Q(\alu_add_sub[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30984_ (.D(_02621_),
    .Q(\alu_add_sub[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30985_ (.D(_02622_),
    .Q(\alu_add_sub[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30986_ (.D(_02592_),
    .Q(\alu_add_sub[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30987_ (.D(_02593_),
    .Q(\alu_add_sub[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30988_ (.D(_02594_),
    .Q(\alu_add_sub[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30989_ (.D(_02595_),
    .Q(\alu_add_sub[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30990_ (.D(_02596_),
    .Q(\alu_add_sub[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30991_ (.D(_02597_),
    .Q(\alu_add_sub[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30992_ (.D(_02598_),
    .Q(\alu_add_sub[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30993_ (.D(_02599_),
    .Q(\alu_add_sub[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30994_ (.D(_02600_),
    .Q(\alu_add_sub[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30995_ (.D(_02601_),
    .Q(\alu_add_sub[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30996_ (.D(_02603_),
    .Q(\alu_add_sub[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30997_ (.D(_02604_),
    .Q(\alu_add_sub[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30998_ (.D(_02605_),
    .Q(\alu_add_sub[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _30999_ (.D(_02606_),
    .Q(\alu_add_sub[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31000_ (.D(_02607_),
    .Q(\alu_add_sub[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31001_ (.D(_02608_),
    .Q(\alu_add_sub[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31002_ (.D(_02609_),
    .Q(\alu_add_sub[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31003_ (.D(_02610_),
    .Q(\alu_add_sub[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31004_ (.D(_02611_),
    .Q(\alu_add_sub[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31005_ (.D(_02612_),
    .Q(\alu_add_sub[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31006_ (.D(_02614_),
    .Q(\alu_add_sub[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31007_ (.D(_02615_),
    .Q(\alu_add_sub[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31008_ (.D(_15246_),
    .Q(\alu_shl[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31009_ (.D(_15247_),
    .Q(\alu_shl[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31010_ (.D(_15248_),
    .Q(\alu_shl[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31011_ (.D(_15249_),
    .Q(\alu_shl[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31012_ (.D(_15250_),
    .Q(\alu_shl[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31013_ (.D(_15251_),
    .Q(\alu_shl[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31014_ (.D(_15252_),
    .Q(\alu_shl[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31015_ (.D(_15253_),
    .Q(\alu_shl[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31016_ (.D(_15254_),
    .Q(\alu_shl[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31017_ (.D(_15255_),
    .Q(\alu_shl[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31018_ (.D(_15256_),
    .Q(\alu_shl[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31019_ (.D(_15257_),
    .Q(\alu_shl[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31020_ (.D(_15258_),
    .Q(\alu_shl[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31021_ (.D(_15259_),
    .Q(\alu_shl[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31022_ (.D(_15260_),
    .Q(\alu_shl[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31023_ (.D(_15261_),
    .Q(\alu_shl[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31024_ (.D(_15262_),
    .Q(\alu_shr[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31025_ (.D(_15273_),
    .Q(\alu_shr[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31026_ (.D(_15284_),
    .Q(\alu_shr[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31027_ (.D(_15287_),
    .Q(\alu_shr[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31028_ (.D(_15288_),
    .Q(\alu_shr[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31029_ (.D(_15289_),
    .Q(\alu_shr[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31030_ (.D(_15290_),
    .Q(\alu_shr[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31031_ (.D(_15291_),
    .Q(\alu_shr[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31032_ (.D(_15292_),
    .Q(\alu_shr[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31033_ (.D(_15293_),
    .Q(\alu_shr[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31034_ (.D(_15263_),
    .Q(\alu_shr[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31035_ (.D(_15264_),
    .Q(\alu_shr[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31036_ (.D(_15265_),
    .Q(\alu_shr[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31037_ (.D(_15266_),
    .Q(\alu_shr[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31038_ (.D(_15267_),
    .Q(\alu_shr[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31039_ (.D(_15268_),
    .Q(\alu_shr[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31040_ (.D(_15269_),
    .Q(\alu_shr[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31041_ (.D(_15270_),
    .Q(\alu_shr[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31042_ (.D(_15271_),
    .Q(\alu_shr[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31043_ (.D(_15272_),
    .Q(\alu_shr[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31044_ (.D(_15274_),
    .Q(\alu_shr[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31045_ (.D(_15275_),
    .Q(\alu_shr[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31046_ (.D(_15276_),
    .Q(\alu_shr[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31047_ (.D(_15277_),
    .Q(\alu_shr[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31048_ (.D(_15278_),
    .Q(\alu_shr[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31049_ (.D(_15279_),
    .Q(\alu_shr[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31050_ (.D(_15280_),
    .Q(\alu_shr[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31051_ (.D(_15281_),
    .Q(\alu_shr[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31052_ (.D(_15282_),
    .Q(\alu_shr[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31053_ (.D(_15283_),
    .Q(\alu_shr[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31054_ (.D(_15285_),
    .Q(\alu_shr[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31055_ (.D(_15286_),
    .Q(\alu_shr[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31056_ (.D(_00000_),
    .Q(alu_eq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31057_ (.D(_00002_),
    .Q(alu_ltu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31058_ (.D(_00001_),
    .Q(alu_lts),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31059_ (.D(_02623_),
    .Q(\pcpi_mul.rd[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31060_ (.D(_02624_),
    .Q(\pcpi_mul.rd[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31061_ (.D(_02625_),
    .Q(\pcpi_mul.rd[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31062_ (.D(_02626_),
    .Q(\pcpi_mul.rd[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31063_ (.D(_02627_),
    .Q(\pcpi_mul.rd[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31064_ (.D(_02628_),
    .Q(\pcpi_mul.rd[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31065_ (.D(_02683_),
    .Q(\pcpi_mul.rd[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31066_ (.D(_02684_),
    .Q(\pcpi_mul.rd[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31067_ (.D(_02685_),
    .Q(\pcpi_mul.rd[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31068_ (.D(_02686_),
    .Q(\pcpi_mul.rd[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31069_ (.D(_02629_),
    .Q(\pcpi_mul.rd[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31070_ (.D(_02630_),
    .Q(\pcpi_mul.rd[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31071_ (.D(_02631_),
    .Q(\pcpi_mul.rd[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31072_ (.D(_02632_),
    .Q(\pcpi_mul.rd[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31073_ (.D(_02633_),
    .Q(\pcpi_mul.rd[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31074_ (.D(_02634_),
    .Q(\pcpi_mul.rd[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31075_ (.D(_02635_),
    .Q(\pcpi_mul.rd[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31076_ (.D(_02636_),
    .Q(\pcpi_mul.rd[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31077_ (.D(_02637_),
    .Q(\pcpi_mul.rd[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31078_ (.D(_02638_),
    .Q(\pcpi_mul.rd[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31079_ (.D(_02639_),
    .Q(\pcpi_mul.rd[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31080_ (.D(_02640_),
    .Q(\pcpi_mul.rd[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31081_ (.D(_02641_),
    .Q(\pcpi_mul.rd[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31082_ (.D(_02642_),
    .Q(\pcpi_mul.rd[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31083_ (.D(_02643_),
    .Q(\pcpi_mul.rd[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31084_ (.D(_02644_),
    .Q(\pcpi_mul.rd[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31085_ (.D(_02645_),
    .Q(\pcpi_mul.rd[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31086_ (.D(_02646_),
    .Q(\pcpi_mul.rd[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31087_ (.D(_02647_),
    .Q(\pcpi_mul.rd[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31088_ (.D(_02648_),
    .Q(\pcpi_mul.rd[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31089_ (.D(_02649_),
    .Q(\pcpi_mul.rd[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31090_ (.D(_02650_),
    .Q(\pcpi_mul.rd[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31091_ (.D(_02651_),
    .Q(\pcpi_mul.rd[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31092_ (.D(_02652_),
    .Q(\pcpi_mul.rd[33] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31093_ (.D(_02653_),
    .Q(\pcpi_mul.rd[34] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31094_ (.D(_02654_),
    .Q(\pcpi_mul.rd[35] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31095_ (.D(_02655_),
    .Q(\pcpi_mul.rd[36] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31096_ (.D(_02656_),
    .Q(\pcpi_mul.rd[37] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31097_ (.D(_02657_),
    .Q(\pcpi_mul.rd[38] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31098_ (.D(_02658_),
    .Q(\pcpi_mul.rd[39] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31099_ (.D(_02659_),
    .Q(\pcpi_mul.rd[40] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31100_ (.D(_02660_),
    .Q(\pcpi_mul.rd[41] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31101_ (.D(_02661_),
    .Q(\pcpi_mul.rd[42] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31102_ (.D(_02662_),
    .Q(\pcpi_mul.rd[43] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31103_ (.D(_02663_),
    .Q(\pcpi_mul.rd[44] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31104_ (.D(_02664_),
    .Q(\pcpi_mul.rd[45] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31105_ (.D(_02665_),
    .Q(\pcpi_mul.rd[46] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31106_ (.D(_02666_),
    .Q(\pcpi_mul.rd[47] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31107_ (.D(_02667_),
    .Q(\pcpi_mul.rd[48] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31108_ (.D(_02668_),
    .Q(\pcpi_mul.rd[49] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31109_ (.D(_02669_),
    .Q(\pcpi_mul.rd[50] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31110_ (.D(_02670_),
    .Q(\pcpi_mul.rd[51] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31111_ (.D(_02671_),
    .Q(\pcpi_mul.rd[52] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31112_ (.D(_02672_),
    .Q(\pcpi_mul.rd[53] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31113_ (.D(_02673_),
    .Q(\pcpi_mul.rd[54] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31114_ (.D(_02674_),
    .Q(\pcpi_mul.rd[55] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31115_ (.D(_02675_),
    .Q(\pcpi_mul.rd[56] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31116_ (.D(_02676_),
    .Q(\pcpi_mul.rd[57] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31117_ (.D(_02677_),
    .Q(\pcpi_mul.rd[58] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31118_ (.D(_02678_),
    .Q(\pcpi_mul.rd[59] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31119_ (.D(_02679_),
    .Q(\pcpi_mul.rd[60] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31120_ (.D(_02680_),
    .Q(\pcpi_mul.rd[61] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31121_ (.D(_02681_),
    .Q(\pcpi_mul.rd[62] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31122_ (.D(_02682_),
    .Q(\pcpi_mul.rd[63] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31123_ (.D(\pcpi_mul.instr_any_mulh ),
    .Q(\pcpi_mul.shift_out ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31124_ (.D(_00038_),
    .Q(\cpu_state[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31125_ (.D(_00039_),
    .Q(\cpu_state[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31126_ (.D(_00040_),
    .Q(\cpu_state[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31127_ (.D(_00041_),
    .Q(\cpu_state[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31128_ (.D(_00042_),
    .Q(\cpu_state[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31129_ (.D(_00043_),
    .Q(\cpu_state[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31130_ (.D(_00044_),
    .Q(\cpu_state[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31131_ (.D(_02771_),
    .Q(\cpuregs[8][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31132_ (.D(_02772_),
    .Q(\cpuregs[8][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31133_ (.D(_02773_),
    .Q(\cpuregs[8][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31134_ (.D(_02774_),
    .Q(\cpuregs[8][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31135_ (.D(_02775_),
    .Q(\cpuregs[8][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31136_ (.D(_02776_),
    .Q(\cpuregs[8][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31137_ (.D(_02777_),
    .Q(\cpuregs[8][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31138_ (.D(_02778_),
    .Q(\cpuregs[8][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31139_ (.D(_02779_),
    .Q(\cpuregs[8][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31140_ (.D(_02780_),
    .Q(\cpuregs[8][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31141_ (.D(_02781_),
    .Q(\cpuregs[8][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31142_ (.D(_02782_),
    .Q(\cpuregs[8][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31143_ (.D(_02783_),
    .Q(\cpuregs[8][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31144_ (.D(_02784_),
    .Q(\cpuregs[8][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31145_ (.D(_02785_),
    .Q(\cpuregs[8][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31146_ (.D(_02786_),
    .Q(\cpuregs[8][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31147_ (.D(_02787_),
    .Q(\cpuregs[8][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31148_ (.D(_02788_),
    .Q(\cpuregs[8][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31149_ (.D(_02789_),
    .Q(\cpuregs[8][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31150_ (.D(_02790_),
    .Q(\cpuregs[8][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31151_ (.D(_02791_),
    .Q(\cpuregs[8][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31152_ (.D(_02792_),
    .Q(\cpuregs[8][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31153_ (.D(_02793_),
    .Q(\cpuregs[8][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31154_ (.D(_02794_),
    .Q(\cpuregs[8][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31155_ (.D(_02795_),
    .Q(\cpuregs[8][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31156_ (.D(_02796_),
    .Q(\cpuregs[8][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31157_ (.D(_02797_),
    .Q(\cpuregs[8][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31158_ (.D(_02798_),
    .Q(\cpuregs[8][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31159_ (.D(_02799_),
    .Q(\cpuregs[8][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31160_ (.D(_02800_),
    .Q(\cpuregs[8][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31161_ (.D(_02801_),
    .Q(\cpuregs[8][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31162_ (.D(_02802_),
    .Q(\cpuregs[8][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31163_ (.D(_02803_),
    .Q(\cpuregs[14][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31164_ (.D(_02804_),
    .Q(\cpuregs[14][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31165_ (.D(_02805_),
    .Q(\cpuregs[14][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31166_ (.D(_02806_),
    .Q(\cpuregs[14][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31167_ (.D(_02807_),
    .Q(\cpuregs[14][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31168_ (.D(_02808_),
    .Q(\cpuregs[14][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31169_ (.D(_02809_),
    .Q(\cpuregs[14][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31170_ (.D(_02810_),
    .Q(\cpuregs[14][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31171_ (.D(_02811_),
    .Q(\cpuregs[14][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31172_ (.D(_02812_),
    .Q(\cpuregs[14][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31173_ (.D(_02813_),
    .Q(\cpuregs[14][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31174_ (.D(_02814_),
    .Q(\cpuregs[14][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31175_ (.D(_02815_),
    .Q(\cpuregs[14][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31176_ (.D(_02816_),
    .Q(\cpuregs[14][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31177_ (.D(_02817_),
    .Q(\cpuregs[14][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31178_ (.D(_02818_),
    .Q(\cpuregs[14][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31179_ (.D(_02819_),
    .Q(\cpuregs[14][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31180_ (.D(_02820_),
    .Q(\cpuregs[14][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31181_ (.D(_02821_),
    .Q(\cpuregs[14][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31182_ (.D(_02822_),
    .Q(\cpuregs[14][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31183_ (.D(_02823_),
    .Q(\cpuregs[14][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31184_ (.D(_02824_),
    .Q(\cpuregs[14][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31185_ (.D(_02825_),
    .Q(\cpuregs[14][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31186_ (.D(_02826_),
    .Q(\cpuregs[14][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31187_ (.D(_02827_),
    .Q(\cpuregs[14][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31188_ (.D(_02828_),
    .Q(\cpuregs[14][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31189_ (.D(_02829_),
    .Q(\cpuregs[14][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31190_ (.D(_02830_),
    .Q(\cpuregs[14][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31191_ (.D(_02831_),
    .Q(\cpuregs[14][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31192_ (.D(_02832_),
    .Q(\cpuregs[14][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31193_ (.D(_02833_),
    .Q(\cpuregs[14][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31194_ (.D(_02834_),
    .Q(\cpuregs[14][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31195_ (.D(_02835_),
    .Q(\cpuregs[0][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31196_ (.D(_02836_),
    .Q(\cpuregs[0][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31197_ (.D(_02837_),
    .Q(\cpuregs[0][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31198_ (.D(_02838_),
    .Q(\cpuregs[0][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31199_ (.D(_02839_),
    .Q(\cpuregs[0][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31200_ (.D(_02840_),
    .Q(\cpuregs[0][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31201_ (.D(_02841_),
    .Q(\cpuregs[0][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31202_ (.D(_02842_),
    .Q(\cpuregs[0][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31203_ (.D(_02843_),
    .Q(\cpuregs[0][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31204_ (.D(_02844_),
    .Q(\cpuregs[0][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31205_ (.D(_02845_),
    .Q(\cpuregs[0][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31206_ (.D(_02846_),
    .Q(\cpuregs[0][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31207_ (.D(_02847_),
    .Q(\cpuregs[0][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31208_ (.D(_02848_),
    .Q(\cpuregs[0][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31209_ (.D(_02849_),
    .Q(\cpuregs[0][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31210_ (.D(_02850_),
    .Q(\cpuregs[0][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31211_ (.D(_02851_),
    .Q(\cpuregs[0][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31212_ (.D(_02852_),
    .Q(\cpuregs[0][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31213_ (.D(_02853_),
    .Q(\cpuregs[0][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31214_ (.D(_02854_),
    .Q(\cpuregs[0][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31215_ (.D(_02855_),
    .Q(\cpuregs[0][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31216_ (.D(_02856_),
    .Q(\cpuregs[0][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31217_ (.D(_02857_),
    .Q(\cpuregs[0][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31218_ (.D(_02858_),
    .Q(\cpuregs[0][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31219_ (.D(_02859_),
    .Q(\cpuregs[0][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31220_ (.D(_02860_),
    .Q(\cpuregs[0][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31221_ (.D(_02861_),
    .Q(\cpuregs[0][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31222_ (.D(_02862_),
    .Q(\cpuregs[0][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31223_ (.D(_02863_),
    .Q(\cpuregs[0][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31224_ (.D(_02864_),
    .Q(\cpuregs[0][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31225_ (.D(_02865_),
    .Q(\cpuregs[0][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31226_ (.D(_02866_),
    .Q(\cpuregs[0][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31227_ (.D(_02867_),
    .Q(\cpuregs[10][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31228_ (.D(_02868_),
    .Q(\cpuregs[10][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31229_ (.D(_02869_),
    .Q(\cpuregs[10][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31230_ (.D(_02870_),
    .Q(\cpuregs[10][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31231_ (.D(_02871_),
    .Q(\cpuregs[10][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31232_ (.D(_02872_),
    .Q(\cpuregs[10][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31233_ (.D(_02873_),
    .Q(\cpuregs[10][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31234_ (.D(_02874_),
    .Q(\cpuregs[10][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31235_ (.D(_02875_),
    .Q(\cpuregs[10][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31236_ (.D(_02876_),
    .Q(\cpuregs[10][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31237_ (.D(_02877_),
    .Q(\cpuregs[10][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31238_ (.D(_02878_),
    .Q(\cpuregs[10][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31239_ (.D(_02879_),
    .Q(\cpuregs[10][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31240_ (.D(_02880_),
    .Q(\cpuregs[10][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31241_ (.D(_02881_),
    .Q(\cpuregs[10][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31242_ (.D(_02882_),
    .Q(\cpuregs[10][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31243_ (.D(_02883_),
    .Q(\cpuregs[10][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31244_ (.D(_02884_),
    .Q(\cpuregs[10][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31245_ (.D(_02885_),
    .Q(\cpuregs[10][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31246_ (.D(_02886_),
    .Q(\cpuregs[10][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31247_ (.D(_02887_),
    .Q(\cpuregs[10][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31248_ (.D(_02888_),
    .Q(\cpuregs[10][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31249_ (.D(_02889_),
    .Q(\cpuregs[10][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31250_ (.D(_02890_),
    .Q(\cpuregs[10][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31251_ (.D(_02891_),
    .Q(\cpuregs[10][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31252_ (.D(_02892_),
    .Q(\cpuregs[10][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31253_ (.D(_02893_),
    .Q(\cpuregs[10][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31254_ (.D(_02894_),
    .Q(\cpuregs[10][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31255_ (.D(_02895_),
    .Q(\cpuregs[10][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31256_ (.D(_02896_),
    .Q(\cpuregs[10][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31257_ (.D(_02897_),
    .Q(\cpuregs[10][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31258_ (.D(_02898_),
    .Q(\cpuregs[10][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31259_ (.D(_02899_),
    .Q(\cpuregs[18][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31260_ (.D(_02900_),
    .Q(\cpuregs[18][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31261_ (.D(_02901_),
    .Q(\cpuregs[18][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31262_ (.D(_02902_),
    .Q(\cpuregs[18][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31263_ (.D(_02903_),
    .Q(\cpuregs[18][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31264_ (.D(_02904_),
    .Q(\cpuregs[18][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31265_ (.D(_02905_),
    .Q(\cpuregs[18][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31266_ (.D(_02906_),
    .Q(\cpuregs[18][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31267_ (.D(_02907_),
    .Q(\cpuregs[18][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31268_ (.D(_02908_),
    .Q(\cpuregs[18][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31269_ (.D(_02909_),
    .Q(\cpuregs[18][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31270_ (.D(_02910_),
    .Q(\cpuregs[18][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31271_ (.D(_02911_),
    .Q(\cpuregs[18][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31272_ (.D(_02912_),
    .Q(\cpuregs[18][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31273_ (.D(_02913_),
    .Q(\cpuregs[18][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31274_ (.D(_02914_),
    .Q(\cpuregs[18][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31275_ (.D(_02915_),
    .Q(\cpuregs[18][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31276_ (.D(_02916_),
    .Q(\cpuregs[18][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31277_ (.D(_02917_),
    .Q(\cpuregs[18][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31278_ (.D(_02918_),
    .Q(\cpuregs[18][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31279_ (.D(_02919_),
    .Q(\cpuregs[18][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31280_ (.D(_02920_),
    .Q(\cpuregs[18][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31281_ (.D(_02921_),
    .Q(\cpuregs[18][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31282_ (.D(_02922_),
    .Q(\cpuregs[18][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31283_ (.D(_02923_),
    .Q(\cpuregs[18][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31284_ (.D(_02924_),
    .Q(\cpuregs[18][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31285_ (.D(_02925_),
    .Q(\cpuregs[18][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31286_ (.D(_02926_),
    .Q(\cpuregs[18][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31287_ (.D(_02927_),
    .Q(\cpuregs[18][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31288_ (.D(_02928_),
    .Q(\cpuregs[18][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31289_ (.D(_02929_),
    .Q(\cpuregs[18][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31290_ (.D(_02930_),
    .Q(\cpuregs[18][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31291_ (.D(_02931_),
    .Q(\mem_rdata_q[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31292_ (.D(_02932_),
    .Q(\mem_rdata_q[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31293_ (.D(_02933_),
    .Q(\mem_rdata_q[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31294_ (.D(_02934_),
    .Q(\mem_rdata_q[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31295_ (.D(_02935_),
    .Q(\mem_rdata_q[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31296_ (.D(_02936_),
    .Q(\mem_rdata_q[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31297_ (.D(_02937_),
    .Q(\mem_rdata_q[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31298_ (.D(_02938_),
    .Q(\mem_rdata_q[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31299_ (.D(_02939_),
    .Q(\mem_rdata_q[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31300_ (.D(_02940_),
    .Q(\mem_rdata_q[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31301_ (.D(_02941_),
    .Q(\mem_rdata_q[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31302_ (.D(_02942_),
    .Q(\mem_rdata_q[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31303_ (.D(_02943_),
    .Q(\mem_rdata_q[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31304_ (.D(_02944_),
    .Q(\mem_rdata_q[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31305_ (.D(_02945_),
    .Q(\mem_rdata_q[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31306_ (.D(_02946_),
    .Q(\mem_rdata_q[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31307_ (.D(_02947_),
    .Q(\mem_rdata_q[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31308_ (.D(_02948_),
    .Q(\mem_rdata_q[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31309_ (.D(_02949_),
    .Q(\mem_rdata_q[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31310_ (.D(_02950_),
    .Q(\mem_rdata_q[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31311_ (.D(_02951_),
    .Q(\mem_rdata_q[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31312_ (.D(_02952_),
    .Q(\mem_rdata_q[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31313_ (.D(_02953_),
    .Q(\mem_rdata_q[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31314_ (.D(_02954_),
    .Q(\mem_rdata_q[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31315_ (.D(_02955_),
    .Q(\mem_rdata_q[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31316_ (.D(_02956_),
    .Q(\mem_rdata_q[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31317_ (.D(_02957_),
    .Q(\mem_rdata_q[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31318_ (.D(_02958_),
    .Q(\mem_rdata_q[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31319_ (.D(_02959_),
    .Q(\mem_rdata_q[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31320_ (.D(_02960_),
    .Q(\mem_rdata_q[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31321_ (.D(_02961_),
    .Q(\mem_rdata_q[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31322_ (.D(_02962_),
    .Q(\mem_rdata_q[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31323_ (.D(_02963_),
    .Q(\cpuregs[2][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31324_ (.D(_02964_),
    .Q(\cpuregs[2][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31325_ (.D(_02965_),
    .Q(\cpuregs[2][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31326_ (.D(_02966_),
    .Q(\cpuregs[2][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31327_ (.D(_02967_),
    .Q(\cpuregs[2][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31328_ (.D(_02968_),
    .Q(\cpuregs[2][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31329_ (.D(_02969_),
    .Q(\cpuregs[2][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31330_ (.D(_02970_),
    .Q(\cpuregs[2][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31331_ (.D(_02971_),
    .Q(\cpuregs[2][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31332_ (.D(_02972_),
    .Q(\cpuregs[2][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31333_ (.D(_02973_),
    .Q(\cpuregs[2][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31334_ (.D(_02974_),
    .Q(\cpuregs[2][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31335_ (.D(_02975_),
    .Q(\cpuregs[2][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31336_ (.D(_02976_),
    .Q(\cpuregs[2][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31337_ (.D(_02977_),
    .Q(\cpuregs[2][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31338_ (.D(_02978_),
    .Q(\cpuregs[2][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31339_ (.D(_02979_),
    .Q(\cpuregs[2][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31340_ (.D(_02980_),
    .Q(\cpuregs[2][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31341_ (.D(_02981_),
    .Q(\cpuregs[2][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31342_ (.D(_02982_),
    .Q(\cpuregs[2][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31343_ (.D(_02983_),
    .Q(\cpuregs[2][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31344_ (.D(_02984_),
    .Q(\cpuregs[2][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31345_ (.D(_02985_),
    .Q(\cpuregs[2][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31346_ (.D(_02986_),
    .Q(\cpuregs[2][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31347_ (.D(_02987_),
    .Q(\cpuregs[2][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31348_ (.D(_02988_),
    .Q(\cpuregs[2][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31349_ (.D(_02989_),
    .Q(\cpuregs[2][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31350_ (.D(_02990_),
    .Q(\cpuregs[2][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31351_ (.D(_02991_),
    .Q(\cpuregs[2][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31352_ (.D(_02992_),
    .Q(\cpuregs[2][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31353_ (.D(_02993_),
    .Q(\cpuregs[2][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31354_ (.D(_02994_),
    .Q(\cpuregs[2][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31355_ (.D(_02995_),
    .Q(\cpuregs[5][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31356_ (.D(_02996_),
    .Q(\cpuregs[5][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31357_ (.D(_02997_),
    .Q(\cpuregs[5][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31358_ (.D(_02998_),
    .Q(\cpuregs[5][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31359_ (.D(_02999_),
    .Q(\cpuregs[5][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31360_ (.D(_03000_),
    .Q(\cpuregs[5][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31361_ (.D(_03001_),
    .Q(\cpuregs[5][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31362_ (.D(_03002_),
    .Q(\cpuregs[5][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31363_ (.D(_03003_),
    .Q(\cpuregs[5][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31364_ (.D(_03004_),
    .Q(\cpuregs[5][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31365_ (.D(_03005_),
    .Q(\cpuregs[5][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31366_ (.D(_03006_),
    .Q(\cpuregs[5][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31367_ (.D(_03007_),
    .Q(\cpuregs[5][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31368_ (.D(_03008_),
    .Q(\cpuregs[5][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31369_ (.D(_03009_),
    .Q(\cpuregs[5][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31370_ (.D(_03010_),
    .Q(\cpuregs[5][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31371_ (.D(_03011_),
    .Q(\cpuregs[5][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31372_ (.D(_03012_),
    .Q(\cpuregs[5][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31373_ (.D(_03013_),
    .Q(\cpuregs[5][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31374_ (.D(_03014_),
    .Q(\cpuregs[5][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31375_ (.D(_03015_),
    .Q(\cpuregs[5][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31376_ (.D(_03016_),
    .Q(\cpuregs[5][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31377_ (.D(_03017_),
    .Q(\cpuregs[5][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31378_ (.D(_03018_),
    .Q(\cpuregs[5][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31379_ (.D(_03019_),
    .Q(\cpuregs[5][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31380_ (.D(_03020_),
    .Q(\cpuregs[5][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31381_ (.D(_03021_),
    .Q(\cpuregs[5][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31382_ (.D(_03022_),
    .Q(\cpuregs[5][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31383_ (.D(_03023_),
    .Q(\cpuregs[5][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31384_ (.D(_03024_),
    .Q(\cpuregs[5][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31385_ (.D(_03025_),
    .Q(\cpuregs[5][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31386_ (.D(_03026_),
    .Q(\cpuregs[5][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31387_ (.D(_03027_),
    .Q(\pcpi_mul.rs1[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31388_ (.D(_03028_),
    .Q(\pcpi_mul.rs1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31389_ (.D(_03029_),
    .Q(\pcpi_mul.rs1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31390_ (.D(_03030_),
    .Q(\pcpi_mul.rs1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31391_ (.D(_03031_),
    .Q(\pcpi_mul.rs1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31392_ (.D(_03032_),
    .Q(\pcpi_mul.rs1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31393_ (.D(_03033_),
    .Q(\pcpi_mul.rs1[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31394_ (.D(_03034_),
    .Q(\pcpi_mul.rs1[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31395_ (.D(_03035_),
    .Q(\pcpi_mul.rs1[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31396_ (.D(_03036_),
    .Q(\pcpi_mul.rs1[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31397_ (.D(_03037_),
    .Q(\pcpi_mul.rs1[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31398_ (.D(_03038_),
    .Q(\pcpi_mul.rs1[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31399_ (.D(_03039_),
    .Q(\pcpi_mul.rs1[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31400_ (.D(_03040_),
    .Q(\pcpi_mul.rs1[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31401_ (.D(_03041_),
    .Q(\pcpi_mul.rs1[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31402_ (.D(_03042_),
    .Q(\pcpi_mul.rs1[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31403_ (.D(_03043_),
    .Q(\pcpi_mul.rs1[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31404_ (.D(_03044_),
    .Q(\pcpi_mul.rs1[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31405_ (.D(_03045_),
    .Q(\pcpi_mul.rs1[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31406_ (.D(_03046_),
    .Q(\pcpi_mul.rs1[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31407_ (.D(_03047_),
    .Q(\pcpi_mul.rs1[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31408_ (.D(_03048_),
    .Q(\pcpi_mul.rs1[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31409_ (.D(_03049_),
    .Q(\pcpi_mul.rs1[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31410_ (.D(_03050_),
    .Q(\pcpi_mul.rs1[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31411_ (.D(_03051_),
    .Q(\pcpi_mul.rs1[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31412_ (.D(_03052_),
    .Q(\pcpi_mul.rs1[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31413_ (.D(_03053_),
    .Q(\pcpi_mul.rs1[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31414_ (.D(_03054_),
    .Q(\pcpi_mul.rs1[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31415_ (.D(_03055_),
    .Q(\pcpi_mul.rs1[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31416_ (.D(_03056_),
    .Q(\pcpi_mul.rs1[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31417_ (.D(_03057_),
    .Q(\pcpi_mul.rs1[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31418_ (.D(_03058_),
    .Q(\pcpi_mul.rs1[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31419_ (.D(_03059_),
    .Q(net156),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31420_ (.D(_03060_),
    .Q(net159),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31421_ (.D(_03061_),
    .Q(net160),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31422_ (.D(_03062_),
    .Q(net161),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31423_ (.D(_03063_),
    .Q(net162),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31424_ (.D(_03064_),
    .Q(net163),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31425_ (.D(_03065_),
    .Q(net164),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31426_ (.D(_03066_),
    .Q(net165),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31427_ (.D(_03067_),
    .Q(net135),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31428_ (.D(_03068_),
    .Q(net136),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31429_ (.D(_03069_),
    .Q(net137),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31430_ (.D(_03070_),
    .Q(net138),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31431_ (.D(_03071_),
    .Q(net139),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31432_ (.D(_03072_),
    .Q(net140),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31433_ (.D(_03073_),
    .Q(net141),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31434_ (.D(_03074_),
    .Q(net142),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31435_ (.D(_03075_),
    .Q(net143),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31436_ (.D(_03076_),
    .Q(net144),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31437_ (.D(_03077_),
    .Q(net146),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31438_ (.D(_03078_),
    .Q(net147),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31439_ (.D(_03079_),
    .Q(net148),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31440_ (.D(_03080_),
    .Q(net149),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31441_ (.D(_03081_),
    .Q(net150),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31442_ (.D(_03082_),
    .Q(net151),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31443_ (.D(_03083_),
    .Q(net152),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31444_ (.D(_03084_),
    .Q(net153),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31445_ (.D(_03085_),
    .Q(net154),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31446_ (.D(_03086_),
    .Q(net155),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31447_ (.D(_03087_),
    .Q(net157),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31448_ (.D(_03088_),
    .Q(net158),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31449_ (.D(_03089_),
    .Q(net306),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31450_ (.D(_03090_),
    .Q(net317),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31451_ (.D(_03091_),
    .Q(net328),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31452_ (.D(_03092_),
    .Q(net331),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31453_ (.D(_03093_),
    .Q(net332),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31454_ (.D(_03094_),
    .Q(net333),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31455_ (.D(_03095_),
    .Q(net334),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31456_ (.D(_03096_),
    .Q(net335),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31457_ (.D(_03097_),
    .Q(net336),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31458_ (.D(_03098_),
    .Q(net337),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31459_ (.D(_03099_),
    .Q(net307),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31460_ (.D(_03100_),
    .Q(net308),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31461_ (.D(_03101_),
    .Q(net309),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31462_ (.D(_03102_),
    .Q(net310),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31463_ (.D(_03103_),
    .Q(net311),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31464_ (.D(_03104_),
    .Q(net312),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31465_ (.D(_03105_),
    .Q(net313),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31466_ (.D(_03106_),
    .Q(net314),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31467_ (.D(_03107_),
    .Q(net315),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31468_ (.D(_03108_),
    .Q(net316),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31469_ (.D(_03109_),
    .Q(net318),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31470_ (.D(_03110_),
    .Q(net319),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31471_ (.D(_03111_),
    .Q(net320),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31472_ (.D(_03112_),
    .Q(net321),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31473_ (.D(_03113_),
    .Q(net322),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31474_ (.D(_03114_),
    .Q(net323),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31475_ (.D(_03115_),
    .Q(net324),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31476_ (.D(_03116_),
    .Q(net325),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31477_ (.D(_03117_),
    .Q(net326),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31478_ (.D(_03118_),
    .Q(net327),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31479_ (.D(_03119_),
    .Q(net329),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31480_ (.D(_03120_),
    .Q(net330),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31481_ (.D(_03121_),
    .Q(net274),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31482_ (.D(_03122_),
    .Q(net285),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31483_ (.D(_03123_),
    .Q(net296),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31484_ (.D(_03124_),
    .Q(net299),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31485_ (.D(_03125_),
    .Q(net300),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31486_ (.D(_03126_),
    .Q(net301),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31487_ (.D(_03127_),
    .Q(net302),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31488_ (.D(_03128_),
    .Q(net303),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31489_ (.D(_03129_),
    .Q(net304),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31490_ (.D(_03130_),
    .Q(net305),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31491_ (.D(_03131_),
    .Q(net275),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31492_ (.D(_03132_),
    .Q(net276),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31493_ (.D(_03133_),
    .Q(net277),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31494_ (.D(_03134_),
    .Q(net278),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31495_ (.D(_03135_),
    .Q(net279),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31496_ (.D(_03136_),
    .Q(net280),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31497_ (.D(_03137_),
    .Q(net281),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31498_ (.D(_03138_),
    .Q(net282),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31499_ (.D(_03139_),
    .Q(net283),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31500_ (.D(_03140_),
    .Q(net284),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31501_ (.D(_03141_),
    .Q(net286),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31502_ (.D(_03142_),
    .Q(net287),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31503_ (.D(_03143_),
    .Q(net288),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31504_ (.D(_03144_),
    .Q(net289),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31505_ (.D(_03145_),
    .Q(net290),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31506_ (.D(_03146_),
    .Q(net291),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31507_ (.D(_03147_),
    .Q(net292),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31508_ (.D(_03148_),
    .Q(net293),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31509_ (.D(_03149_),
    .Q(net294),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31510_ (.D(_03150_),
    .Q(net295),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31511_ (.D(_03151_),
    .Q(net297),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31512_ (.D(_03152_),
    .Q(net298),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31513_ (.D(_03153_),
    .Q(instr_lui),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31514_ (.D(_03154_),
    .Q(instr_auipc),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31515_ (.D(_03155_),
    .Q(instr_jal),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31516_ (.D(_03156_),
    .Q(instr_jalr),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31517_ (.D(_03157_),
    .Q(instr_lb),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31518_ (.D(_03158_),
    .Q(instr_lh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31519_ (.D(_03159_),
    .Q(instr_lw),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31520_ (.D(_03160_),
    .Q(instr_lbu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31521_ (.D(_03161_),
    .Q(instr_lhu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31522_ (.D(_03162_),
    .Q(instr_sb),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31523_ (.D(_03163_),
    .Q(instr_sh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31524_ (.D(_03164_),
    .Q(instr_sw),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31525_ (.D(_03165_),
    .Q(instr_slli),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31526_ (.D(_03166_),
    .Q(instr_srli),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31527_ (.D(_03167_),
    .Q(instr_srai),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31528_ (.D(_03168_),
    .Q(instr_rdcycle),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31529_ (.D(_03169_),
    .Q(instr_rdcycleh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31530_ (.D(_03170_),
    .Q(instr_rdinstr),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31531_ (.D(_03171_),
    .Q(instr_rdinstrh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31532_ (.D(_03172_),
    .Q(instr_ecall_ebreak),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31533_ (.D(_03173_),
    .Q(instr_getq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31534_ (.D(_03174_),
    .Q(instr_setq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31535_ (.D(_03175_),
    .Q(instr_retirq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31536_ (.D(_03176_),
    .Q(instr_maskirq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31537_ (.D(_03177_),
    .Q(instr_waitirq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31538_ (.D(_03178_),
    .Q(instr_timer),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31539_ (.D(_03179_),
    .Q(\decoded_rd[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31540_ (.D(_03180_),
    .Q(\decoded_rd[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31541_ (.D(_03181_),
    .Q(\decoded_rd[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31542_ (.D(_03182_),
    .Q(\decoded_rd[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31543_ (.D(_03183_),
    .Q(\decoded_rd[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31544_ (.D(_03184_),
    .Q(\decoded_imm[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31545_ (.D(_03185_),
    .Q(\decoded_imm_uj[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31546_ (.D(_03186_),
    .Q(\decoded_imm_uj[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31547_ (.D(_03187_),
    .Q(\decoded_imm_uj[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31548_ (.D(_03188_),
    .Q(\decoded_imm_uj[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31549_ (.D(_03189_),
    .Q(\decoded_imm_uj[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31550_ (.D(_03190_),
    .Q(\decoded_imm_uj[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31551_ (.D(_03191_),
    .Q(\decoded_imm_uj[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31552_ (.D(_03192_),
    .Q(\decoded_imm_uj[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31553_ (.D(_03193_),
    .Q(\decoded_imm_uj[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31554_ (.D(_03194_),
    .Q(\decoded_imm_uj[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31555_ (.D(_03195_),
    .Q(\decoded_imm_uj[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31556_ (.D(_03196_),
    .Q(\decoded_imm_uj[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31557_ (.D(_03197_),
    .Q(\decoded_imm_uj[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31558_ (.D(_03198_),
    .Q(\decoded_imm_uj[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31559_ (.D(_03199_),
    .Q(\decoded_imm_uj[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31560_ (.D(_03200_),
    .Q(\decoded_imm_uj[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31561_ (.D(_03201_),
    .Q(\decoded_imm_uj[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31562_ (.D(_03202_),
    .Q(\decoded_imm_uj[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31563_ (.D(_03203_),
    .Q(\decoded_imm_uj[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31564_ (.D(_03204_),
    .Q(\decoded_imm_uj[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31565_ (.D(_03205_),
    .Q(is_lb_lh_lw_lbu_lhu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31566_ (.D(_03206_),
    .Q(is_slli_srli_srai),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31567_ (.D(_03207_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31568_ (.D(_03208_),
    .Q(is_sb_sh_sw),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31569_ (.D(_03209_),
    .Q(\cpuregs[13][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31570_ (.D(_03210_),
    .Q(\cpuregs[13][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31571_ (.D(_03211_),
    .Q(\cpuregs[13][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31572_ (.D(_03212_),
    .Q(\cpuregs[13][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31573_ (.D(_03213_),
    .Q(\cpuregs[13][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31574_ (.D(_03214_),
    .Q(\cpuregs[13][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31575_ (.D(_03215_),
    .Q(\cpuregs[13][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31576_ (.D(_03216_),
    .Q(\cpuregs[13][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31577_ (.D(_03217_),
    .Q(\cpuregs[13][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31578_ (.D(_03218_),
    .Q(\cpuregs[13][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31579_ (.D(_03219_),
    .Q(\cpuregs[13][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31580_ (.D(_03220_),
    .Q(\cpuregs[13][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31581_ (.D(_03221_),
    .Q(\cpuregs[13][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31582_ (.D(_03222_),
    .Q(\cpuregs[13][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31583_ (.D(_03223_),
    .Q(\cpuregs[13][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31584_ (.D(_03224_),
    .Q(\cpuregs[13][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31585_ (.D(_03225_),
    .Q(\cpuregs[13][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31586_ (.D(_03226_),
    .Q(\cpuregs[13][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31587_ (.D(_03227_),
    .Q(\cpuregs[13][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31588_ (.D(_03228_),
    .Q(\cpuregs[13][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31589_ (.D(_03229_),
    .Q(\cpuregs[13][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31590_ (.D(_03230_),
    .Q(\cpuregs[13][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31591_ (.D(_03231_),
    .Q(\cpuregs[13][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31592_ (.D(_03232_),
    .Q(\cpuregs[13][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31593_ (.D(_03233_),
    .Q(\cpuregs[13][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31594_ (.D(_03234_),
    .Q(\cpuregs[13][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31595_ (.D(_03235_),
    .Q(\cpuregs[13][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31596_ (.D(_03236_),
    .Q(\cpuregs[13][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31597_ (.D(_03237_),
    .Q(\cpuregs[13][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31598_ (.D(_03238_),
    .Q(\cpuregs[13][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31599_ (.D(_03239_),
    .Q(\cpuregs[13][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31600_ (.D(_03240_),
    .Q(\cpuregs[13][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31601_ (.D(_03241_),
    .Q(is_alu_reg_imm),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31602_ (.D(_03242_),
    .Q(is_alu_reg_reg),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31603_ (.D(_03243_),
    .Q(net270),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31604_ (.D(_03244_),
    .Q(net271),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31605_ (.D(_03245_),
    .Q(net272),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31606_ (.D(_03246_),
    .Q(net273),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31607_ (.D(_03247_),
    .Q(\pcpi_mul.rs2[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31608_ (.D(_03248_),
    .Q(\pcpi_mul.rs2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31609_ (.D(_03249_),
    .Q(\pcpi_mul.rs2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31610_ (.D(_03250_),
    .Q(\pcpi_mul.rs2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31611_ (.D(_03251_),
    .Q(\pcpi_mul.rs2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31612_ (.D(_03252_),
    .Q(\pcpi_mul.rs2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31613_ (.D(_03253_),
    .Q(\pcpi_mul.rs2[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31614_ (.D(_03254_),
    .Q(\pcpi_mul.rs2[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31615_ (.D(_03255_),
    .Q(\pcpi_mul.rs2[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31616_ (.D(_03256_),
    .Q(\pcpi_mul.rs2[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31617_ (.D(_03257_),
    .Q(\pcpi_mul.rs2[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31618_ (.D(_03258_),
    .Q(\pcpi_mul.rs2[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31619_ (.D(_03259_),
    .Q(\pcpi_mul.rs2[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31620_ (.D(_03260_),
    .Q(\pcpi_mul.rs2[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31621_ (.D(_03261_),
    .Q(\pcpi_mul.rs2[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31622_ (.D(_03262_),
    .Q(\pcpi_mul.rs2[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31623_ (.D(_03263_),
    .Q(\pcpi_mul.rs2[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31624_ (.D(_03264_),
    .Q(\pcpi_mul.rs2[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31625_ (.D(_03265_),
    .Q(\pcpi_mul.rs2[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31626_ (.D(_03266_),
    .Q(\pcpi_mul.rs2[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31627_ (.D(_03267_),
    .Q(\pcpi_mul.rs2[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31628_ (.D(_03268_),
    .Q(\pcpi_mul.rs2[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31629_ (.D(_03269_),
    .Q(\pcpi_mul.rs2[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31630_ (.D(_03270_),
    .Q(\pcpi_mul.rs2[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31631_ (.D(_03271_),
    .Q(\pcpi_mul.rs2[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31632_ (.D(_03272_),
    .Q(\pcpi_mul.rs2[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31633_ (.D(_03273_),
    .Q(\pcpi_mul.rs2[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31634_ (.D(_03274_),
    .Q(\pcpi_mul.rs2[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31635_ (.D(_03275_),
    .Q(\pcpi_mul.rs2[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31636_ (.D(_03276_),
    .Q(\pcpi_mul.rs2[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31637_ (.D(_03277_),
    .Q(\pcpi_mul.rs2[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31638_ (.D(_03278_),
    .Q(\pcpi_mul.rs2[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31639_ (.D(_03279_),
    .Q(\cpuregs[17][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31640_ (.D(_03280_),
    .Q(\cpuregs[17][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31641_ (.D(_03281_),
    .Q(\cpuregs[17][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31642_ (.D(_03282_),
    .Q(\cpuregs[17][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31643_ (.D(_03283_),
    .Q(\cpuregs[17][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31644_ (.D(_03284_),
    .Q(\cpuregs[17][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31645_ (.D(_03285_),
    .Q(\cpuregs[17][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31646_ (.D(_03286_),
    .Q(\cpuregs[17][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31647_ (.D(_03287_),
    .Q(\cpuregs[17][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31648_ (.D(_03288_),
    .Q(\cpuregs[17][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31649_ (.D(_03289_),
    .Q(\cpuregs[17][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31650_ (.D(_03290_),
    .Q(\cpuregs[17][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31651_ (.D(_03291_),
    .Q(\cpuregs[17][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31652_ (.D(_03292_),
    .Q(\cpuregs[17][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31653_ (.D(_03293_),
    .Q(\cpuregs[17][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31654_ (.D(_03294_),
    .Q(\cpuregs[17][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31655_ (.D(_03295_),
    .Q(\cpuregs[17][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31656_ (.D(_03296_),
    .Q(\cpuregs[17][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31657_ (.D(_03297_),
    .Q(\cpuregs[17][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31658_ (.D(_03298_),
    .Q(\cpuregs[17][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31659_ (.D(_03299_),
    .Q(\cpuregs[17][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31660_ (.D(_03300_),
    .Q(\cpuregs[17][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31661_ (.D(_03301_),
    .Q(\cpuregs[17][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31662_ (.D(_03302_),
    .Q(\cpuregs[17][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31663_ (.D(_03303_),
    .Q(\cpuregs[17][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31664_ (.D(_03304_),
    .Q(\cpuregs[17][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31665_ (.D(_03305_),
    .Q(\cpuregs[17][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31666_ (.D(_03306_),
    .Q(\cpuregs[17][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31667_ (.D(_03307_),
    .Q(\cpuregs[17][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31668_ (.D(_03308_),
    .Q(\cpuregs[17][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31669_ (.D(_03309_),
    .Q(\cpuregs[17][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31670_ (.D(_03310_),
    .Q(\cpuregs[17][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31671_ (.D(_03311_),
    .Q(\cpuregs[16][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31672_ (.D(_03312_),
    .Q(\cpuregs[16][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31673_ (.D(_03313_),
    .Q(\cpuregs[16][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31674_ (.D(_03314_),
    .Q(\cpuregs[16][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31675_ (.D(_03315_),
    .Q(\cpuregs[16][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31676_ (.D(_03316_),
    .Q(\cpuregs[16][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31677_ (.D(_03317_),
    .Q(\cpuregs[16][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31678_ (.D(_03318_),
    .Q(\cpuregs[16][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31679_ (.D(_03319_),
    .Q(\cpuregs[16][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31680_ (.D(_03320_),
    .Q(\cpuregs[16][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31681_ (.D(_03321_),
    .Q(\cpuregs[16][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31682_ (.D(_03322_),
    .Q(\cpuregs[16][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31683_ (.D(_03323_),
    .Q(\cpuregs[16][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31684_ (.D(_03324_),
    .Q(\cpuregs[16][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31685_ (.D(_03325_),
    .Q(\cpuregs[16][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31686_ (.D(_03326_),
    .Q(\cpuregs[16][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31687_ (.D(_03327_),
    .Q(\cpuregs[16][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31688_ (.D(_03328_),
    .Q(\cpuregs[16][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31689_ (.D(_03329_),
    .Q(\cpuregs[16][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31690_ (.D(_03330_),
    .Q(\cpuregs[16][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31691_ (.D(_03331_),
    .Q(\cpuregs[16][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31692_ (.D(_03332_),
    .Q(\cpuregs[16][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31693_ (.D(_03333_),
    .Q(\cpuregs[16][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31694_ (.D(_03334_),
    .Q(\cpuregs[16][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31695_ (.D(_03335_),
    .Q(\cpuregs[16][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31696_ (.D(_03336_),
    .Q(\cpuregs[16][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31697_ (.D(_03337_),
    .Q(\cpuregs[16][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31698_ (.D(_03338_),
    .Q(\cpuregs[16][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31699_ (.D(_03339_),
    .Q(\cpuregs[16][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31700_ (.D(_03340_),
    .Q(\cpuregs[16][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31701_ (.D(_03341_),
    .Q(\cpuregs[16][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31702_ (.D(_03342_),
    .Q(\cpuregs[16][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31703_ (.D(_03343_),
    .Q(\cpuregs[12][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31704_ (.D(_03344_),
    .Q(\cpuregs[12][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31705_ (.D(_03345_),
    .Q(\cpuregs[12][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31706_ (.D(_03346_),
    .Q(\cpuregs[12][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31707_ (.D(_03347_),
    .Q(\cpuregs[12][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31708_ (.D(_03348_),
    .Q(\cpuregs[12][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31709_ (.D(_03349_),
    .Q(\cpuregs[12][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31710_ (.D(_03350_),
    .Q(\cpuregs[12][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31711_ (.D(_03351_),
    .Q(\cpuregs[12][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31712_ (.D(_03352_),
    .Q(\cpuregs[12][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31713_ (.D(_03353_),
    .Q(\cpuregs[12][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31714_ (.D(_03354_),
    .Q(\cpuregs[12][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31715_ (.D(_03355_),
    .Q(\cpuregs[12][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31716_ (.D(_03356_),
    .Q(\cpuregs[12][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31717_ (.D(_03357_),
    .Q(\cpuregs[12][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31718_ (.D(_03358_),
    .Q(\cpuregs[12][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31719_ (.D(_03359_),
    .Q(\cpuregs[12][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31720_ (.D(_03360_),
    .Q(\cpuregs[12][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31721_ (.D(_03361_),
    .Q(\cpuregs[12][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31722_ (.D(_03362_),
    .Q(\cpuregs[12][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31723_ (.D(_03363_),
    .Q(\cpuregs[12][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31724_ (.D(_03364_),
    .Q(\cpuregs[12][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31725_ (.D(_03365_),
    .Q(\cpuregs[12][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31726_ (.D(_03366_),
    .Q(\cpuregs[12][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31727_ (.D(_03367_),
    .Q(\cpuregs[12][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31728_ (.D(_03368_),
    .Q(\cpuregs[12][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31729_ (.D(_03369_),
    .Q(\cpuregs[12][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31730_ (.D(_03370_),
    .Q(\cpuregs[12][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31731_ (.D(_03371_),
    .Q(\cpuregs[12][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31732_ (.D(_03372_),
    .Q(\cpuregs[12][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31733_ (.D(_03373_),
    .Q(\cpuregs[12][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31734_ (.D(_03374_),
    .Q(\cpuregs[12][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31735_ (.D(_03375_),
    .Q(\cpuregs[1][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31736_ (.D(_03376_),
    .Q(\cpuregs[1][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31737_ (.D(_03377_),
    .Q(\cpuregs[1][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31738_ (.D(_03378_),
    .Q(\cpuregs[1][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31739_ (.D(_03379_),
    .Q(\cpuregs[1][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31740_ (.D(_03380_),
    .Q(\cpuregs[1][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31741_ (.D(_03381_),
    .Q(\cpuregs[1][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31742_ (.D(_03382_),
    .Q(\cpuregs[1][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31743_ (.D(_03383_),
    .Q(\cpuregs[1][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31744_ (.D(_03384_),
    .Q(\cpuregs[1][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31745_ (.D(_03385_),
    .Q(\cpuregs[1][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31746_ (.D(_03386_),
    .Q(\cpuregs[1][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31747_ (.D(_03387_),
    .Q(\cpuregs[1][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31748_ (.D(_03388_),
    .Q(\cpuregs[1][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31749_ (.D(_03389_),
    .Q(\cpuregs[1][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31750_ (.D(_03390_),
    .Q(\cpuregs[1][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31751_ (.D(_03391_),
    .Q(\cpuregs[1][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31752_ (.D(_03392_),
    .Q(\cpuregs[1][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31753_ (.D(_03393_),
    .Q(\cpuregs[1][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31754_ (.D(_03394_),
    .Q(\cpuregs[1][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31755_ (.D(_03395_),
    .Q(\cpuregs[1][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31756_ (.D(_03396_),
    .Q(\cpuregs[1][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31757_ (.D(_03397_),
    .Q(\cpuregs[1][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31758_ (.D(_03398_),
    .Q(\cpuregs[1][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31759_ (.D(_03399_),
    .Q(\cpuregs[1][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31760_ (.D(_03400_),
    .Q(\cpuregs[1][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31761_ (.D(_03401_),
    .Q(\cpuregs[1][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31762_ (.D(_03402_),
    .Q(\cpuregs[1][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31763_ (.D(_03403_),
    .Q(\cpuregs[1][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31764_ (.D(_03404_),
    .Q(\cpuregs[1][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31765_ (.D(_03405_),
    .Q(\cpuregs[1][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31766_ (.D(_03406_),
    .Q(\cpuregs[1][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31767_ (.D(_03407_),
    .Q(\cpuregs[3][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31768_ (.D(_03408_),
    .Q(\cpuregs[3][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31769_ (.D(_03409_),
    .Q(\cpuregs[3][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31770_ (.D(_03410_),
    .Q(\cpuregs[3][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31771_ (.D(_03411_),
    .Q(\cpuregs[3][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31772_ (.D(_03412_),
    .Q(\cpuregs[3][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31773_ (.D(_03413_),
    .Q(\cpuregs[3][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31774_ (.D(_03414_),
    .Q(\cpuregs[3][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31775_ (.D(_03415_),
    .Q(\cpuregs[3][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31776_ (.D(_03416_),
    .Q(\cpuregs[3][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31777_ (.D(_03417_),
    .Q(\cpuregs[3][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31778_ (.D(_03418_),
    .Q(\cpuregs[3][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31779_ (.D(_03419_),
    .Q(\cpuregs[3][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31780_ (.D(_03420_),
    .Q(\cpuregs[3][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31781_ (.D(_03421_),
    .Q(\cpuregs[3][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31782_ (.D(_03422_),
    .Q(\cpuregs[3][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31783_ (.D(_03423_),
    .Q(\cpuregs[3][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31784_ (.D(_03424_),
    .Q(\cpuregs[3][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31785_ (.D(_03425_),
    .Q(\cpuregs[3][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31786_ (.D(_03426_),
    .Q(\cpuregs[3][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31787_ (.D(_03427_),
    .Q(\cpuregs[3][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31788_ (.D(_03428_),
    .Q(\cpuregs[3][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31789_ (.D(_03429_),
    .Q(\cpuregs[3][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31790_ (.D(_03430_),
    .Q(\cpuregs[3][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31791_ (.D(_03431_),
    .Q(\cpuregs[3][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31792_ (.D(_03432_),
    .Q(\cpuregs[3][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31793_ (.D(_03433_),
    .Q(\cpuregs[3][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31794_ (.D(_03434_),
    .Q(\cpuregs[3][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31795_ (.D(_03435_),
    .Q(\cpuregs[3][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31796_ (.D(_03436_),
    .Q(\cpuregs[3][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31797_ (.D(_03437_),
    .Q(\cpuregs[3][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31798_ (.D(_03438_),
    .Q(\cpuregs[3][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31799_ (.D(_03439_),
    .Q(\cpuregs[11][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31800_ (.D(_03440_),
    .Q(\cpuregs[11][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31801_ (.D(_03441_),
    .Q(\cpuregs[11][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31802_ (.D(_03442_),
    .Q(\cpuregs[11][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31803_ (.D(_03443_),
    .Q(\cpuregs[11][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31804_ (.D(_03444_),
    .Q(\cpuregs[11][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31805_ (.D(_03445_),
    .Q(\cpuregs[11][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31806_ (.D(_03446_),
    .Q(\cpuregs[11][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31807_ (.D(_03447_),
    .Q(\cpuregs[11][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31808_ (.D(_03448_),
    .Q(\cpuregs[11][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31809_ (.D(_03449_),
    .Q(\cpuregs[11][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31810_ (.D(_03450_),
    .Q(\cpuregs[11][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31811_ (.D(_03451_),
    .Q(\cpuregs[11][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31812_ (.D(_03452_),
    .Q(\cpuregs[11][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31813_ (.D(_03453_),
    .Q(\cpuregs[11][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31814_ (.D(_03454_),
    .Q(\cpuregs[11][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31815_ (.D(_03455_),
    .Q(\cpuregs[11][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31816_ (.D(_03456_),
    .Q(\cpuregs[11][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31817_ (.D(_03457_),
    .Q(\cpuregs[11][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31818_ (.D(_03458_),
    .Q(\cpuregs[11][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31819_ (.D(_03459_),
    .Q(\cpuregs[11][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31820_ (.D(_03460_),
    .Q(\cpuregs[11][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31821_ (.D(_03461_),
    .Q(\cpuregs[11][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31822_ (.D(_03462_),
    .Q(\cpuregs[11][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31823_ (.D(_03463_),
    .Q(\cpuregs[11][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31824_ (.D(_03464_),
    .Q(\cpuregs[11][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31825_ (.D(_03465_),
    .Q(\cpuregs[11][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31826_ (.D(_03466_),
    .Q(\cpuregs[11][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31827_ (.D(_03467_),
    .Q(\cpuregs[11][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31828_ (.D(_03468_),
    .Q(\cpuregs[11][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31829_ (.D(_03469_),
    .Q(\cpuregs[11][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31830_ (.D(_03470_),
    .Q(\cpuregs[11][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31831_ (.D(_03471_),
    .Q(\cpuregs[15][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31832_ (.D(_03472_),
    .Q(\cpuregs[15][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31833_ (.D(_03473_),
    .Q(\cpuregs[15][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31834_ (.D(_03474_),
    .Q(\cpuregs[15][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31835_ (.D(_03475_),
    .Q(\cpuregs[15][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31836_ (.D(_03476_),
    .Q(\cpuregs[15][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31837_ (.D(_03477_),
    .Q(\cpuregs[15][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31838_ (.D(_03478_),
    .Q(\cpuregs[15][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31839_ (.D(_03479_),
    .Q(\cpuregs[15][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31840_ (.D(_03480_),
    .Q(\cpuregs[15][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31841_ (.D(_03481_),
    .Q(\cpuregs[15][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31842_ (.D(_03482_),
    .Q(\cpuregs[15][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31843_ (.D(_03483_),
    .Q(\cpuregs[15][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31844_ (.D(_03484_),
    .Q(\cpuregs[15][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31845_ (.D(_03485_),
    .Q(\cpuregs[15][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31846_ (.D(_03486_),
    .Q(\cpuregs[15][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31847_ (.D(_03487_),
    .Q(\cpuregs[15][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31848_ (.D(_03488_),
    .Q(\cpuregs[15][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31849_ (.D(_03489_),
    .Q(\cpuregs[15][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31850_ (.D(_03490_),
    .Q(\cpuregs[15][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31851_ (.D(_03491_),
    .Q(\cpuregs[15][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31852_ (.D(_03492_),
    .Q(\cpuregs[15][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31853_ (.D(_03493_),
    .Q(\cpuregs[15][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31854_ (.D(_03494_),
    .Q(\cpuregs[15][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31855_ (.D(_03495_),
    .Q(\cpuregs[15][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31856_ (.D(_03496_),
    .Q(\cpuregs[15][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31857_ (.D(_03497_),
    .Q(\cpuregs[15][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31858_ (.D(_03498_),
    .Q(\cpuregs[15][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31859_ (.D(_03499_),
    .Q(\cpuregs[15][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31860_ (.D(_03500_),
    .Q(\cpuregs[15][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31861_ (.D(_03501_),
    .Q(\cpuregs[15][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31862_ (.D(_03502_),
    .Q(\cpuregs[15][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31863_ (.D(_03503_),
    .Q(\latched_rd[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31864_ (.D(_03504_),
    .Q(\cpuregs[7][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31865_ (.D(_03505_),
    .Q(\cpuregs[7][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31866_ (.D(_03506_),
    .Q(\cpuregs[7][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31867_ (.D(_03507_),
    .Q(\cpuregs[7][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31868_ (.D(_03508_),
    .Q(\cpuregs[7][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31869_ (.D(_03509_),
    .Q(\cpuregs[7][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31870_ (.D(_03510_),
    .Q(\cpuregs[7][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31871_ (.D(_03511_),
    .Q(\cpuregs[7][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31872_ (.D(_03512_),
    .Q(\cpuregs[7][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31873_ (.D(_03513_),
    .Q(\cpuregs[7][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31874_ (.D(_03514_),
    .Q(\cpuregs[7][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31875_ (.D(_03515_),
    .Q(\cpuregs[7][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31876_ (.D(_03516_),
    .Q(\cpuregs[7][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31877_ (.D(_03517_),
    .Q(\cpuregs[7][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31878_ (.D(_03518_),
    .Q(\cpuregs[7][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31879_ (.D(_03519_),
    .Q(\cpuregs[7][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31880_ (.D(_03520_),
    .Q(\cpuregs[7][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31881_ (.D(_03521_),
    .Q(\cpuregs[7][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31882_ (.D(_03522_),
    .Q(\cpuregs[7][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31883_ (.D(_03523_),
    .Q(\cpuregs[7][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31884_ (.D(_03524_),
    .Q(\cpuregs[7][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31885_ (.D(_03525_),
    .Q(\cpuregs[7][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31886_ (.D(_03526_),
    .Q(\cpuregs[7][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31887_ (.D(_03527_),
    .Q(\cpuregs[7][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31888_ (.D(_03528_),
    .Q(\cpuregs[7][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31889_ (.D(_03529_),
    .Q(\cpuregs[7][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31890_ (.D(_03530_),
    .Q(\cpuregs[7][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31891_ (.D(_03531_),
    .Q(\cpuregs[7][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31892_ (.D(_03532_),
    .Q(\cpuregs[7][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31893_ (.D(_03533_),
    .Q(\cpuregs[7][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31894_ (.D(_03534_),
    .Q(\cpuregs[7][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31895_ (.D(_03535_),
    .Q(\cpuregs[7][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31896_ (.D(_03536_),
    .Q(net238),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31897_ (.D(_03537_),
    .Q(net249),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31898_ (.D(_03538_),
    .Q(net260),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31899_ (.D(_03539_),
    .Q(net263),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31900_ (.D(_03540_),
    .Q(net264),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31901_ (.D(_03541_),
    .Q(net265),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31902_ (.D(_03542_),
    .Q(net266),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31903_ (.D(_03543_),
    .Q(net267),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31904_ (.D(_03544_),
    .Q(net268),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31905_ (.D(_03545_),
    .Q(net269),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31906_ (.D(_03546_),
    .Q(net239),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31907_ (.D(_03547_),
    .Q(net240),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31908_ (.D(_03548_),
    .Q(net241),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31909_ (.D(_03549_),
    .Q(net242),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31910_ (.D(_03550_),
    .Q(net243),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31911_ (.D(_03551_),
    .Q(net244),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31912_ (.D(_03552_),
    .Q(net245),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31913_ (.D(_03553_),
    .Q(net246),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31914_ (.D(_03554_),
    .Q(net247),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31915_ (.D(_03555_),
    .Q(net248),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31916_ (.D(_03556_),
    .Q(net250),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31917_ (.D(_03557_),
    .Q(net251),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31918_ (.D(_03558_),
    .Q(net252),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31919_ (.D(_03559_),
    .Q(net253),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31920_ (.D(_03560_),
    .Q(net254),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31921_ (.D(_03561_),
    .Q(net255),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31922_ (.D(_03562_),
    .Q(net256),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31923_ (.D(_03563_),
    .Q(net257),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _31924_ (.D(_03564_),
    .Q(net258),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31925_ (.D(_03565_),
    .Q(net259),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31926_ (.D(_03566_),
    .Q(net261),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31927_ (.D(_03567_),
    .Q(net262),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31928_ (.D(_03568_),
    .Q(\cpuregs[19][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31929_ (.D(_03569_),
    .Q(\cpuregs[19][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31930_ (.D(_03570_),
    .Q(\cpuregs[19][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31931_ (.D(_03571_),
    .Q(\cpuregs[19][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31932_ (.D(_03572_),
    .Q(\cpuregs[19][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31933_ (.D(_03573_),
    .Q(\cpuregs[19][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31934_ (.D(_03574_),
    .Q(\cpuregs[19][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31935_ (.D(_03575_),
    .Q(\cpuregs[19][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31936_ (.D(_03576_),
    .Q(\cpuregs[19][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31937_ (.D(_03577_),
    .Q(\cpuregs[19][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31938_ (.D(_03578_),
    .Q(\cpuregs[19][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31939_ (.D(_03579_),
    .Q(\cpuregs[19][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31940_ (.D(_03580_),
    .Q(\cpuregs[19][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31941_ (.D(_03581_),
    .Q(\cpuregs[19][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31942_ (.D(_03582_),
    .Q(\cpuregs[19][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31943_ (.D(_03583_),
    .Q(\cpuregs[19][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31944_ (.D(_03584_),
    .Q(\cpuregs[19][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31945_ (.D(_03585_),
    .Q(\cpuregs[19][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31946_ (.D(_03586_),
    .Q(\cpuregs[19][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31947_ (.D(_03587_),
    .Q(\cpuregs[19][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31948_ (.D(_03588_),
    .Q(\cpuregs[19][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31949_ (.D(_03589_),
    .Q(\cpuregs[19][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31950_ (.D(_03590_),
    .Q(\cpuregs[19][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31951_ (.D(_03591_),
    .Q(\cpuregs[19][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31952_ (.D(_03592_),
    .Q(\cpuregs[19][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31953_ (.D(_03593_),
    .Q(\cpuregs[19][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31954_ (.D(_03594_),
    .Q(\cpuregs[19][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31955_ (.D(_03595_),
    .Q(\cpuregs[19][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31956_ (.D(_03596_),
    .Q(\cpuregs[19][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31957_ (.D(_03597_),
    .Q(\cpuregs[19][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31958_ (.D(_03598_),
    .Q(\cpuregs[19][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31959_ (.D(_03599_),
    .Q(\cpuregs[19][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31960_ (.D(_03600_),
    .Q(\cpuregs[4][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31961_ (.D(_03601_),
    .Q(\cpuregs[4][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31962_ (.D(_03602_),
    .Q(\cpuregs[4][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31963_ (.D(_03603_),
    .Q(\cpuregs[4][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31964_ (.D(_03604_),
    .Q(\cpuregs[4][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31965_ (.D(_03605_),
    .Q(\cpuregs[4][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31966_ (.D(_03606_),
    .Q(\cpuregs[4][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31967_ (.D(_03607_),
    .Q(\cpuregs[4][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31968_ (.D(_03608_),
    .Q(\cpuregs[4][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31969_ (.D(_03609_),
    .Q(\cpuregs[4][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31970_ (.D(_03610_),
    .Q(\cpuregs[4][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31971_ (.D(_03611_),
    .Q(\cpuregs[4][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31972_ (.D(_03612_),
    .Q(\cpuregs[4][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31973_ (.D(_03613_),
    .Q(\cpuregs[4][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31974_ (.D(_03614_),
    .Q(\cpuregs[4][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31975_ (.D(_03615_),
    .Q(\cpuregs[4][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31976_ (.D(_03616_),
    .Q(\cpuregs[4][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31977_ (.D(_03617_),
    .Q(\cpuregs[4][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31978_ (.D(_03618_),
    .Q(\cpuregs[4][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31979_ (.D(_03619_),
    .Q(\cpuregs[4][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31980_ (.D(_03620_),
    .Q(\cpuregs[4][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31981_ (.D(_03621_),
    .Q(\cpuregs[4][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31982_ (.D(_03622_),
    .Q(\cpuregs[4][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31983_ (.D(_03623_),
    .Q(\cpuregs[4][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31984_ (.D(_03624_),
    .Q(\cpuregs[4][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31985_ (.D(_03625_),
    .Q(\cpuregs[4][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31986_ (.D(_03626_),
    .Q(\cpuregs[4][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31987_ (.D(_03627_),
    .Q(\cpuregs[4][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31988_ (.D(_03628_),
    .Q(\cpuregs[4][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31989_ (.D(_03629_),
    .Q(\cpuregs[4][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31990_ (.D(_03630_),
    .Q(\cpuregs[4][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _31991_ (.D(_03631_),
    .Q(\cpuregs[4][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31992_ (.D(_03632_),
    .Q(net200),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31993_ (.D(_03633_),
    .Q(net211),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31994_ (.D(_03634_),
    .Q(net222),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31995_ (.D(_03635_),
    .Q(net225),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31996_ (.D(_03636_),
    .Q(net226),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31997_ (.D(_03637_),
    .Q(net227),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31998_ (.D(_03638_),
    .Q(net228),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _31999_ (.D(_03639_),
    .Q(net229),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32000_ (.D(_03640_),
    .Q(net368),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32001_ (.D(_03641_),
    .Q(net369),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32002_ (.D(_03642_),
    .Q(net339),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32003_ (.D(_03643_),
    .Q(net340),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32004_ (.D(_03644_),
    .Q(net341),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32005_ (.D(_03645_),
    .Q(net342),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32006_ (.D(_03646_),
    .Q(net343),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32007_ (.D(_03647_),
    .Q(net344),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32008_ (.D(_03648_),
    .Q(net345),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32009_ (.D(_03649_),
    .Q(net346),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32010_ (.D(_03650_),
    .Q(net347),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32011_ (.D(_03651_),
    .Q(net348),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32012_ (.D(_03652_),
    .Q(net350),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32013_ (.D(_03653_),
    .Q(net351),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32014_ (.D(_03654_),
    .Q(net352),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32015_ (.D(_03655_),
    .Q(net353),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32016_ (.D(_03656_),
    .Q(net354),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32017_ (.D(_03657_),
    .Q(net355),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32018_ (.D(_03658_),
    .Q(net356),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32019_ (.D(_03659_),
    .Q(net357),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32020_ (.D(_03660_),
    .Q(net358),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32021_ (.D(_03661_),
    .Q(net359),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32022_ (.D(_03662_),
    .Q(net361),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32023_ (.D(_03663_),
    .Q(net362),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32024_ (.D(_03664_),
    .Q(\cpuregs[9][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32025_ (.D(_03665_),
    .Q(\cpuregs[9][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32026_ (.D(_03666_),
    .Q(\cpuregs[9][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32027_ (.D(_03667_),
    .Q(\cpuregs[9][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32028_ (.D(_03668_),
    .Q(\cpuregs[9][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32029_ (.D(_03669_),
    .Q(\cpuregs[9][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32030_ (.D(_03670_),
    .Q(\cpuregs[9][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32031_ (.D(_03671_),
    .Q(\cpuregs[9][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32032_ (.D(_03672_),
    .Q(\cpuregs[9][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32033_ (.D(_03673_),
    .Q(\cpuregs[9][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32034_ (.D(_03674_),
    .Q(\cpuregs[9][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32035_ (.D(_03675_),
    .Q(\cpuregs[9][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32036_ (.D(_03676_),
    .Q(\cpuregs[9][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32037_ (.D(_03677_),
    .Q(\cpuregs[9][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32038_ (.D(_03678_),
    .Q(\cpuregs[9][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32039_ (.D(_03679_),
    .Q(\cpuregs[9][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32040_ (.D(_03680_),
    .Q(\cpuregs[9][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32041_ (.D(_03681_),
    .Q(\cpuregs[9][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32042_ (.D(_03682_),
    .Q(\cpuregs[9][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32043_ (.D(_03683_),
    .Q(\cpuregs[9][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32044_ (.D(_03684_),
    .Q(\cpuregs[9][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32045_ (.D(_03685_),
    .Q(\cpuregs[9][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32046_ (.D(_03686_),
    .Q(\cpuregs[9][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32047_ (.D(_03687_),
    .Q(\cpuregs[9][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32048_ (.D(_03688_),
    .Q(\cpuregs[9][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32049_ (.D(_03689_),
    .Q(\cpuregs[9][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32050_ (.D(_03690_),
    .Q(\cpuregs[9][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32051_ (.D(_03691_),
    .Q(\cpuregs[9][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32052_ (.D(_03692_),
    .Q(\cpuregs[9][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32053_ (.D(_03693_),
    .Q(\cpuregs[9][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32054_ (.D(_03694_),
    .Q(\cpuregs[9][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32055_ (.D(_03695_),
    .Q(\cpuregs[9][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32056_ (.D(_03696_),
    .Q(\cpuregs[6][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32057_ (.D(_03697_),
    .Q(\cpuregs[6][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32058_ (.D(_03698_),
    .Q(\cpuregs[6][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32059_ (.D(_03699_),
    .Q(\cpuregs[6][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32060_ (.D(_03700_),
    .Q(\cpuregs[6][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32061_ (.D(_03701_),
    .Q(\cpuregs[6][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32062_ (.D(_03702_),
    .Q(\cpuregs[6][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32063_ (.D(_03703_),
    .Q(\cpuregs[6][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32064_ (.D(_03704_),
    .Q(\cpuregs[6][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32065_ (.D(_03705_),
    .Q(\cpuregs[6][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32066_ (.D(_03706_),
    .Q(\cpuregs[6][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32067_ (.D(_03707_),
    .Q(\cpuregs[6][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32068_ (.D(_03708_),
    .Q(\cpuregs[6][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32069_ (.D(_03709_),
    .Q(\cpuregs[6][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32070_ (.D(_03710_),
    .Q(\cpuregs[6][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32071_ (.D(_03711_),
    .Q(\cpuregs[6][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32072_ (.D(_03712_),
    .Q(\cpuregs[6][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32073_ (.D(_03713_),
    .Q(\cpuregs[6][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32074_ (.D(_03714_),
    .Q(\cpuregs[6][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32075_ (.D(_03715_),
    .Q(\cpuregs[6][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32076_ (.D(_03716_),
    .Q(\cpuregs[6][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32077_ (.D(_03717_),
    .Q(\cpuregs[6][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32078_ (.D(_03718_),
    .Q(\cpuregs[6][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32079_ (.D(_03719_),
    .Q(\cpuregs[6][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32080_ (.D(_03720_),
    .Q(\cpuregs[6][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32081_ (.D(_03721_),
    .Q(\cpuregs[6][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32082_ (.D(_03722_),
    .Q(\cpuregs[6][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32083_ (.D(_03723_),
    .Q(\cpuregs[6][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32084_ (.D(_03724_),
    .Q(\cpuregs[6][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32085_ (.D(_03725_),
    .Q(\cpuregs[6][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32086_ (.D(_03726_),
    .Q(\cpuregs[6][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32087_ (.D(_03727_),
    .Q(\cpuregs[6][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32088_ (.D(_03728_),
    .Q(\pcpi_mul.active[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32089_ (.D(_03729_),
    .Q(\pcpi_mul.active[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32090_ (.D(_03730_),
    .Q(net408),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32091_ (.D(_03731_),
    .Q(\count_cycle[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32092_ (.D(_03732_),
    .Q(\count_cycle[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32093_ (.D(_03733_),
    .Q(\count_cycle[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32094_ (.D(_03734_),
    .Q(\count_cycle[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32095_ (.D(_03735_),
    .Q(\count_cycle[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32096_ (.D(_03736_),
    .Q(\count_cycle[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32097_ (.D(_03737_),
    .Q(\count_cycle[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32098_ (.D(_03738_),
    .Q(\count_cycle[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32099_ (.D(_03739_),
    .Q(\count_cycle[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32100_ (.D(_03740_),
    .Q(\count_cycle[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32101_ (.D(_03741_),
    .Q(\count_cycle[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32102_ (.D(_03742_),
    .Q(\count_cycle[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32103_ (.D(_03743_),
    .Q(\count_cycle[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32104_ (.D(_03744_),
    .Q(\count_cycle[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32105_ (.D(_03745_),
    .Q(\count_cycle[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32106_ (.D(_03746_),
    .Q(\count_cycle[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32107_ (.D(_03747_),
    .Q(\count_cycle[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32108_ (.D(_03748_),
    .Q(\count_cycle[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32109_ (.D(_03749_),
    .Q(\count_cycle[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32110_ (.D(_03750_),
    .Q(\count_cycle[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32111_ (.D(_03751_),
    .Q(\count_cycle[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32112_ (.D(_03752_),
    .Q(\count_cycle[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32113_ (.D(_03753_),
    .Q(\count_cycle[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32114_ (.D(_03754_),
    .Q(\count_cycle[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32115_ (.D(_03755_),
    .Q(\count_cycle[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32116_ (.D(_03756_),
    .Q(\count_cycle[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32117_ (.D(_03757_),
    .Q(\count_cycle[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32118_ (.D(_03758_),
    .Q(\count_cycle[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32119_ (.D(_03759_),
    .Q(\count_cycle[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32120_ (.D(_03760_),
    .Q(\count_cycle[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32121_ (.D(_03761_),
    .Q(\count_cycle[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32122_ (.D(_03762_),
    .Q(\count_cycle[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32123_ (.D(_03763_),
    .Q(\count_cycle[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32124_ (.D(_03764_),
    .Q(\count_cycle[33] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32125_ (.D(_03765_),
    .Q(\count_cycle[34] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32126_ (.D(_03766_),
    .Q(\count_cycle[35] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32127_ (.D(_03767_),
    .Q(\count_cycle[36] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32128_ (.D(_03768_),
    .Q(\count_cycle[37] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32129_ (.D(_03769_),
    .Q(\count_cycle[38] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32130_ (.D(_03770_),
    .Q(\count_cycle[39] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32131_ (.D(_03771_),
    .Q(\count_cycle[40] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32132_ (.D(_03772_),
    .Q(\count_cycle[41] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32133_ (.D(_03773_),
    .Q(\count_cycle[42] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32134_ (.D(_03774_),
    .Q(\count_cycle[43] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32135_ (.D(_03775_),
    .Q(\count_cycle[44] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32136_ (.D(_03776_),
    .Q(\count_cycle[45] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32137_ (.D(_03777_),
    .Q(\count_cycle[46] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32138_ (.D(_03778_),
    .Q(\count_cycle[47] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32139_ (.D(_03779_),
    .Q(\count_cycle[48] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32140_ (.D(_03780_),
    .Q(\count_cycle[49] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32141_ (.D(_03781_),
    .Q(\count_cycle[50] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32142_ (.D(_03782_),
    .Q(\count_cycle[51] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32143_ (.D(_03783_),
    .Q(\count_cycle[52] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32144_ (.D(_03784_),
    .Q(\count_cycle[53] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32145_ (.D(_03785_),
    .Q(\count_cycle[54] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32146_ (.D(_03786_),
    .Q(\count_cycle[55] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32147_ (.D(_03787_),
    .Q(\count_cycle[56] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32148_ (.D(_03788_),
    .Q(\count_cycle[57] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32149_ (.D(_03789_),
    .Q(\count_cycle[58] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32150_ (.D(_03790_),
    .Q(\count_cycle[59] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32151_ (.D(_03791_),
    .Q(\count_cycle[60] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32152_ (.D(_03792_),
    .Q(\count_cycle[61] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32153_ (.D(_03793_),
    .Q(\count_cycle[62] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32154_ (.D(_03794_),
    .Q(\count_cycle[63] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32155_ (.D(_03795_),
    .Q(\timer[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32156_ (.D(_03796_),
    .Q(\timer[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32157_ (.D(_03797_),
    .Q(\timer[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32158_ (.D(_03798_),
    .Q(\timer[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32159_ (.D(_03799_),
    .Q(\timer[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32160_ (.D(_03800_),
    .Q(\timer[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32161_ (.D(_03801_),
    .Q(\timer[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32162_ (.D(_03802_),
    .Q(\timer[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32163_ (.D(_03803_),
    .Q(\timer[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32164_ (.D(_03804_),
    .Q(\timer[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32165_ (.D(_03805_),
    .Q(\timer[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32166_ (.D(_03806_),
    .Q(\timer[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32167_ (.D(_03807_),
    .Q(\timer[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32168_ (.D(_03808_),
    .Q(\timer[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32169_ (.D(_03809_),
    .Q(\timer[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32170_ (.D(_03810_),
    .Q(\timer[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32171_ (.D(_03811_),
    .Q(\timer[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32172_ (.D(_03812_),
    .Q(\timer[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32173_ (.D(_03813_),
    .Q(\timer[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32174_ (.D(_03814_),
    .Q(\timer[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32175_ (.D(_03815_),
    .Q(\timer[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32176_ (.D(_03816_),
    .Q(\timer[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32177_ (.D(_03817_),
    .Q(\timer[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32178_ (.D(_03818_),
    .Q(\timer[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32179_ (.D(_03819_),
    .Q(\timer[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32180_ (.D(_03820_),
    .Q(\timer[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32181_ (.D(_03821_),
    .Q(\timer[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32182_ (.D(_03822_),
    .Q(\timer[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32183_ (.D(_03823_),
    .Q(\timer[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32184_ (.D(_03824_),
    .Q(\timer[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32185_ (.D(_03825_),
    .Q(\timer[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32186_ (.D(_03826_),
    .Q(\timer[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32187_ (.D(_03827_),
    .Q(pcpi_timeout),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32188_ (.D(_03828_),
    .Q(decoder_pseudo_trigger),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32189_ (.D(_03829_),
    .Q(is_compare),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32190_ (.D(_03830_),
    .Q(do_waitirq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32191_ (.D(_03831_),
    .Q(net237),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32192_ (.D(_03832_),
    .Q(net370),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32193_ (.D(_03833_),
    .Q(net102),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32194_ (.D(_03834_),
    .Q(net113),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32195_ (.D(_03835_),
    .Q(net124),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32196_ (.D(_03836_),
    .Q(net127),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32197_ (.D(_03837_),
    .Q(net128),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32198_ (.D(_03838_),
    .Q(net129),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32199_ (.D(_03839_),
    .Q(net130),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32200_ (.D(_03840_),
    .Q(net131),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32201_ (.D(_03841_),
    .Q(net132),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32202_ (.D(_03842_),
    .Q(net133),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32203_ (.D(_03843_),
    .Q(net103),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32204_ (.D(_03844_),
    .Q(net104),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32205_ (.D(_03845_),
    .Q(net105),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32206_ (.D(_03846_),
    .Q(net106),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32207_ (.D(_03847_),
    .Q(net107),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32208_ (.D(_03848_),
    .Q(net108),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32209_ (.D(_03849_),
    .Q(net109),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32210_ (.D(_03850_),
    .Q(net110),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32211_ (.D(_03851_),
    .Q(net111),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32212_ (.D(_03852_),
    .Q(net112),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32213_ (.D(_03853_),
    .Q(net114),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32214_ (.D(_03854_),
    .Q(net115),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32215_ (.D(_03855_),
    .Q(net116),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32216_ (.D(_03856_),
    .Q(net117),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32217_ (.D(_03857_),
    .Q(net118),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32218_ (.D(_03858_),
    .Q(net119),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32219_ (.D(_03859_),
    .Q(net120),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32220_ (.D(_03860_),
    .Q(net121),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32221_ (.D(_03861_),
    .Q(net122),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32222_ (.D(_03862_),
    .Q(net123),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32223_ (.D(_03863_),
    .Q(net125),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32224_ (.D(_03864_),
    .Q(net126),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32225_ (.D(_03865_),
    .Q(\count_instr[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32226_ (.D(_03866_),
    .Q(\count_instr[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32227_ (.D(_03867_),
    .Q(\count_instr[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32228_ (.D(_03868_),
    .Q(\count_instr[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32229_ (.D(_03869_),
    .Q(\count_instr[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32230_ (.D(_03870_),
    .Q(\count_instr[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32231_ (.D(_03871_),
    .Q(\count_instr[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32232_ (.D(_03872_),
    .Q(\count_instr[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32233_ (.D(_03873_),
    .Q(\count_instr[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32234_ (.D(_03874_),
    .Q(\count_instr[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32235_ (.D(_03875_),
    .Q(\count_instr[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32236_ (.D(_03876_),
    .Q(\count_instr[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32237_ (.D(_03877_),
    .Q(\count_instr[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32238_ (.D(_03878_),
    .Q(\count_instr[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32239_ (.D(_03879_),
    .Q(\count_instr[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32240_ (.D(_03880_),
    .Q(\count_instr[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32241_ (.D(_03881_),
    .Q(\count_instr[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32242_ (.D(_03882_),
    .Q(\count_instr[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32243_ (.D(_03883_),
    .Q(\count_instr[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32244_ (.D(_03884_),
    .Q(\count_instr[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32245_ (.D(_03885_),
    .Q(\count_instr[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32246_ (.D(_03886_),
    .Q(\count_instr[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32247_ (.D(_03887_),
    .Q(\count_instr[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32248_ (.D(_03888_),
    .Q(\count_instr[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32249_ (.D(_03889_),
    .Q(\count_instr[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32250_ (.D(_03890_),
    .Q(\count_instr[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32251_ (.D(_03891_),
    .Q(\count_instr[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32252_ (.D(_03892_),
    .Q(\count_instr[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32253_ (.D(_03893_),
    .Q(\count_instr[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32254_ (.D(_03894_),
    .Q(\count_instr[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32255_ (.D(_03895_),
    .Q(\count_instr[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32256_ (.D(_03896_),
    .Q(\count_instr[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32257_ (.D(_03897_),
    .Q(\count_instr[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32258_ (.D(_03898_),
    .Q(\count_instr[33] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32259_ (.D(_03899_),
    .Q(\count_instr[34] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32260_ (.D(_03900_),
    .Q(\count_instr[35] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32261_ (.D(_03901_),
    .Q(\count_instr[36] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32262_ (.D(_03902_),
    .Q(\count_instr[37] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32263_ (.D(_03903_),
    .Q(\count_instr[38] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32264_ (.D(_03904_),
    .Q(\count_instr[39] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32265_ (.D(_03905_),
    .Q(\count_instr[40] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32266_ (.D(_03906_),
    .Q(\count_instr[41] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32267_ (.D(_03907_),
    .Q(\count_instr[42] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32268_ (.D(_03908_),
    .Q(\count_instr[43] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32269_ (.D(_03909_),
    .Q(\count_instr[44] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32270_ (.D(_03910_),
    .Q(\count_instr[45] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32271_ (.D(_03911_),
    .Q(\count_instr[46] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32272_ (.D(_03912_),
    .Q(\count_instr[47] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32273_ (.D(_03913_),
    .Q(\count_instr[48] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32274_ (.D(_03914_),
    .Q(\count_instr[49] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32275_ (.D(_03915_),
    .Q(\count_instr[50] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32276_ (.D(_03916_),
    .Q(\count_instr[51] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32277_ (.D(_03917_),
    .Q(\count_instr[52] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32278_ (.D(_03918_),
    .Q(\count_instr[53] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32279_ (.D(_03919_),
    .Q(\count_instr[54] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32280_ (.D(_03920_),
    .Q(\count_instr[55] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32281_ (.D(_03921_),
    .Q(\count_instr[56] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32282_ (.D(_03922_),
    .Q(\count_instr[57] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32283_ (.D(_03923_),
    .Q(\count_instr[58] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32284_ (.D(_03924_),
    .Q(\count_instr[59] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32285_ (.D(_03925_),
    .Q(\count_instr[60] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32286_ (.D(_03926_),
    .Q(\count_instr[61] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32287_ (.D(_03927_),
    .Q(\count_instr[62] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32288_ (.D(_03928_),
    .Q(\count_instr[63] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32289_ (.D(_03929_),
    .Q(\reg_pc[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32290_ (.D(_03930_),
    .Q(\reg_pc[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32291_ (.D(_03931_),
    .Q(\reg_pc[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32292_ (.D(_03932_),
    .Q(\reg_pc[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32293_ (.D(_03933_),
    .Q(\reg_pc[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32294_ (.D(_03934_),
    .Q(\reg_pc[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32295_ (.D(_03935_),
    .Q(\reg_pc[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32296_ (.D(_03936_),
    .Q(\reg_pc[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32297_ (.D(_03937_),
    .Q(\reg_pc[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32298_ (.D(_03938_),
    .Q(\reg_pc[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32299_ (.D(_03939_),
    .Q(\reg_pc[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32300_ (.D(_03940_),
    .Q(\reg_pc[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32301_ (.D(_03941_),
    .Q(\reg_pc[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32302_ (.D(_03942_),
    .Q(\reg_pc[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32303_ (.D(_03943_),
    .Q(\reg_pc[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32304_ (.D(_03944_),
    .Q(\reg_pc[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32305_ (.D(_03945_),
    .Q(\reg_pc[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32306_ (.D(_03946_),
    .Q(\reg_pc[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32307_ (.D(_03947_),
    .Q(\reg_pc[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32308_ (.D(_03948_),
    .Q(\reg_pc[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32309_ (.D(_03949_),
    .Q(\reg_pc[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32310_ (.D(_03950_),
    .Q(\reg_pc[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32311_ (.D(_03951_),
    .Q(\reg_pc[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32312_ (.D(_03952_),
    .Q(\reg_pc[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32313_ (.D(_03953_),
    .Q(\reg_pc[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32314_ (.D(_03954_),
    .Q(\reg_pc[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32315_ (.D(_03955_),
    .Q(\reg_pc[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32316_ (.D(_03956_),
    .Q(\reg_pc[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32317_ (.D(_03957_),
    .Q(\reg_pc[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32318_ (.D(_03958_),
    .Q(\reg_pc[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32319_ (.D(_03959_),
    .Q(\reg_pc[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32320_ (.D(_03960_),
    .Q(\reg_next_pc[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32321_ (.D(_03961_),
    .Q(\reg_next_pc[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32322_ (.D(_03962_),
    .Q(\reg_next_pc[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32323_ (.D(_03963_),
    .Q(\reg_next_pc[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32324_ (.D(_03964_),
    .Q(\reg_next_pc[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32325_ (.D(_03965_),
    .Q(\reg_next_pc[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32326_ (.D(_03966_),
    .Q(\reg_next_pc[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32327_ (.D(_03967_),
    .Q(\reg_next_pc[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32328_ (.D(_03968_),
    .Q(\reg_next_pc[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32329_ (.D(_03969_),
    .Q(\reg_next_pc[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32330_ (.D(_03970_),
    .Q(\reg_next_pc[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32331_ (.D(_03971_),
    .Q(\reg_next_pc[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32332_ (.D(_03972_),
    .Q(\reg_next_pc[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32333_ (.D(_03973_),
    .Q(\reg_next_pc[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32334_ (.D(_03974_),
    .Q(\reg_next_pc[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32335_ (.D(_03975_),
    .Q(\reg_next_pc[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32336_ (.D(_03976_),
    .Q(\reg_next_pc[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32337_ (.D(_03977_),
    .Q(\reg_next_pc[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32338_ (.D(_03978_),
    .Q(\reg_next_pc[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32339_ (.D(_03979_),
    .Q(\reg_next_pc[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32340_ (.D(_03980_),
    .Q(\reg_next_pc[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32341_ (.D(_03981_),
    .Q(\reg_next_pc[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32342_ (.D(_03982_),
    .Q(\reg_next_pc[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32343_ (.D(_03983_),
    .Q(\reg_next_pc[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32344_ (.D(_03984_),
    .Q(\reg_next_pc[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32345_ (.D(_03985_),
    .Q(\reg_next_pc[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32346_ (.D(_03986_),
    .Q(\reg_next_pc[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32347_ (.D(_03987_),
    .Q(\reg_next_pc[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32348_ (.D(_03988_),
    .Q(\reg_next_pc[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32349_ (.D(_03989_),
    .Q(\reg_next_pc[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32350_ (.D(_03990_),
    .Q(\reg_next_pc[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32351_ (.D(_03991_),
    .Q(mem_do_rdata),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32352_ (.D(_03992_),
    .Q(mem_do_wdata),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32353_ (.D(_03993_),
    .Q(\pcpi_timeout_counter[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32354_ (.D(_03994_),
    .Q(\pcpi_timeout_counter[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32355_ (.D(_03995_),
    .Q(\pcpi_timeout_counter[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32356_ (.D(_03996_),
    .Q(\pcpi_timeout_counter[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32357_ (.D(_03997_),
    .Q(instr_beq),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32358_ (.D(_03998_),
    .Q(instr_bne),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32359_ (.D(_03999_),
    .Q(instr_blt),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32360_ (.D(_04000_),
    .Q(instr_bge),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32361_ (.D(_04001_),
    .Q(instr_bltu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32362_ (.D(_04002_),
    .Q(instr_bgeu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32363_ (.D(_04003_),
    .Q(instr_addi),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32364_ (.D(_04004_),
    .Q(instr_slti),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32365_ (.D(_04005_),
    .Q(instr_sltiu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32366_ (.D(_04006_),
    .Q(instr_xori),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32367_ (.D(_04007_),
    .Q(instr_ori),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32368_ (.D(_04008_),
    .Q(instr_andi),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32369_ (.D(_04009_),
    .Q(instr_add),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32370_ (.D(_04010_),
    .Q(instr_sub),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32371_ (.D(_04011_),
    .Q(instr_sll),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32372_ (.D(_04012_),
    .Q(instr_slt),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32373_ (.D(_04013_),
    .Q(instr_sltu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32374_ (.D(_04014_),
    .Q(instr_xor),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32375_ (.D(_04015_),
    .Q(instr_srl),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32376_ (.D(_04016_),
    .Q(instr_sra),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32377_ (.D(_04017_),
    .Q(instr_or),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32378_ (.D(_04018_),
    .Q(instr_and),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32379_ (.D(_04019_),
    .Q(\decoded_rs1[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32380_ (.D(_04020_),
    .Q(\decoded_rs1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32381_ (.D(_04021_),
    .Q(\decoded_rs1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32382_ (.D(_04022_),
    .Q(\decoded_rs1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32383_ (.D(_04023_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32384_ (.D(_04024_),
    .Q(net166),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32385_ (.D(_04025_),
    .Q(\irq_mask[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32386_ (.D(_04026_),
    .Q(\irq_mask[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32387_ (.D(_04027_),
    .Q(\irq_mask[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32388_ (.D(_04028_),
    .Q(\irq_mask[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32389_ (.D(_04029_),
    .Q(\irq_mask[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32390_ (.D(_04030_),
    .Q(\irq_mask[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32391_ (.D(_04031_),
    .Q(\irq_mask[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32392_ (.D(_04032_),
    .Q(\irq_mask[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32393_ (.D(_04033_),
    .Q(\irq_mask[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32394_ (.D(_04034_),
    .Q(\irq_mask[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32395_ (.D(_04035_),
    .Q(\irq_mask[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32396_ (.D(_04036_),
    .Q(\irq_mask[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32397_ (.D(_04037_),
    .Q(\irq_mask[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32398_ (.D(_04038_),
    .Q(\irq_mask[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32399_ (.D(_04039_),
    .Q(\irq_mask[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32400_ (.D(_04040_),
    .Q(\irq_mask[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32401_ (.D(_04041_),
    .Q(\irq_mask[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32402_ (.D(_04042_),
    .Q(\irq_mask[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32403_ (.D(_04043_),
    .Q(\irq_mask[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32404_ (.D(_04044_),
    .Q(\irq_mask[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32405_ (.D(_04045_),
    .Q(\irq_mask[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32406_ (.D(_04046_),
    .Q(\irq_mask[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32407_ (.D(_04047_),
    .Q(\irq_mask[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32408_ (.D(_04048_),
    .Q(\irq_mask[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32409_ (.D(_04049_),
    .Q(\irq_mask[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32410_ (.D(_04050_),
    .Q(\irq_mask[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32411_ (.D(_04051_),
    .Q(\irq_mask[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32412_ (.D(_04052_),
    .Q(\irq_mask[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32413_ (.D(_04053_),
    .Q(\irq_mask[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32414_ (.D(_04054_),
    .Q(\irq_mask[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32415_ (.D(_04055_),
    .Q(\irq_mask[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32416_ (.D(_04056_),
    .Q(\irq_mask[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32417_ (.D(_04057_),
    .Q(mem_do_prefetch),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32418_ (.D(_04058_),
    .Q(mem_do_rinst),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32419_ (.D(_04059_),
    .Q(\irq_state[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32420_ (.D(_04060_),
    .Q(\irq_state[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32421_ (.D(_04061_),
    .Q(latched_store),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32422_ (.D(_04062_),
    .Q(latched_stalu),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32423_ (.D(_04063_),
    .Q(\pcpi_mul.rs2[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32424_ (.D(_04064_),
    .Q(\pcpi_mul.rs1[32] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32425_ (.D(_04065_),
    .Q(irq_delay),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32426_ (.D(_04066_),
    .Q(\decoded_rs1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32427_ (.D(_04067_),
    .Q(\mem_state[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 _32428_ (.D(_04068_),
    .Q(\mem_state[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32429_ (.D(_04069_),
    .Q(latched_branch),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32430_ (.D(_04070_),
    .Q(latched_is_lh),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _32431_ (.D(_04071_),
    .Q(latched_is_lb),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 _32432_ (.D(_04072_),
    .Q(irq_active),
    .CLK(clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7707 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(irq[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(irq[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(irq[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(irq[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(irq[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(irq[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(irq[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(irq[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(irq[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(irq[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(irq[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(irq[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(irq[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_6 input14 (.A(irq[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(irq[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(irq[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(irq[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(irq[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(irq[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(irq[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(irq[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_6 input22 (.A(irq[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(irq[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(irq[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_8 input25 (.A(irq[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_6 input26 (.A(irq[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(irq[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(irq[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(irq[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(irq[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(irq[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_6 input32 (.A(irq[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(mem_rdata[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(mem_rdata[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_6 input35 (.A(mem_rdata[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_8 input36 (.A(mem_rdata[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(mem_rdata[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_6 input38 (.A(mem_rdata[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(mem_rdata[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_8 input40 (.A(mem_rdata[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(mem_rdata[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_6 input42 (.A(mem_rdata[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(mem_rdata[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_8 input44 (.A(mem_rdata[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_8 input45 (.A(mem_rdata[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(mem_rdata[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_8 input47 (.A(mem_rdata[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_6 input48 (.A(mem_rdata[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_6 input49 (.A(mem_rdata[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_6 input50 (.A(mem_rdata[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_8 input51 (.A(mem_rdata[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_6 input52 (.A(mem_rdata[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_6 input53 (.A(mem_rdata[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_6 input54 (.A(mem_rdata[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_6 input55 (.A(mem_rdata[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(mem_rdata[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(mem_rdata[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_6 input58 (.A(mem_rdata[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_6 input59 (.A(mem_rdata[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_8 input60 (.A(mem_rdata[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 input61 (.A(mem_rdata[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_6 input62 (.A(mem_rdata[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_6 input63 (.A(mem_rdata[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 input64 (.A(mem_rdata[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_8 input65 (.A(mem_ready),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(pcpi_rd[0]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(pcpi_rd[10]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(pcpi_rd[11]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(pcpi_rd[12]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(pcpi_rd[13]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(pcpi_rd[14]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(pcpi_rd[15]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(pcpi_rd[16]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(pcpi_rd[17]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(pcpi_rd[18]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(pcpi_rd[19]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(pcpi_rd[1]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(pcpi_rd[20]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(pcpi_rd[21]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(pcpi_rd[22]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(pcpi_rd[23]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(pcpi_rd[24]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(pcpi_rd[25]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(pcpi_rd[26]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(pcpi_rd[27]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(pcpi_rd[28]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(pcpi_rd[29]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(pcpi_rd[2]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(pcpi_rd[30]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(pcpi_rd[31]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(pcpi_rd[3]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(pcpi_rd[4]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(pcpi_rd[5]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(pcpi_rd[6]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(pcpi_rd[7]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(pcpi_rd[8]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(pcpi_rd[9]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(pcpi_ready),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(pcpi_wait),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(pcpi_wr),
    .X(net100));
 sky130_fd_sc_hd__buf_6 input101 (.A(resetn),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(eoi[0]));
 sky130_fd_sc_hd__clkbuf_2 output103 (.A(net103),
    .X(eoi[10]));
 sky130_fd_sc_hd__clkbuf_2 output104 (.A(net104),
    .X(eoi[11]));
 sky130_fd_sc_hd__clkbuf_2 output105 (.A(net105),
    .X(eoi[12]));
 sky130_fd_sc_hd__clkbuf_2 output106 (.A(net106),
    .X(eoi[13]));
 sky130_fd_sc_hd__clkbuf_2 output107 (.A(net107),
    .X(eoi[14]));
 sky130_fd_sc_hd__clkbuf_2 output108 (.A(net108),
    .X(eoi[15]));
 sky130_fd_sc_hd__clkbuf_2 output109 (.A(net109),
    .X(eoi[16]));
 sky130_fd_sc_hd__clkbuf_2 output110 (.A(net110),
    .X(eoi[17]));
 sky130_fd_sc_hd__clkbuf_2 output111 (.A(net111),
    .X(eoi[18]));
 sky130_fd_sc_hd__clkbuf_2 output112 (.A(net112),
    .X(eoi[19]));
 sky130_fd_sc_hd__clkbuf_2 output113 (.A(net113),
    .X(eoi[1]));
 sky130_fd_sc_hd__clkbuf_2 output114 (.A(net114),
    .X(eoi[20]));
 sky130_fd_sc_hd__clkbuf_2 output115 (.A(net115),
    .X(eoi[21]));
 sky130_fd_sc_hd__clkbuf_2 output116 (.A(net116),
    .X(eoi[22]));
 sky130_fd_sc_hd__clkbuf_2 output117 (.A(net117),
    .X(eoi[23]));
 sky130_fd_sc_hd__clkbuf_2 output118 (.A(net118),
    .X(eoi[24]));
 sky130_fd_sc_hd__clkbuf_2 output119 (.A(net119),
    .X(eoi[25]));
 sky130_fd_sc_hd__clkbuf_2 output120 (.A(net120),
    .X(eoi[26]));
 sky130_fd_sc_hd__clkbuf_2 output121 (.A(net121),
    .X(eoi[27]));
 sky130_fd_sc_hd__clkbuf_2 output122 (.A(net122),
    .X(eoi[28]));
 sky130_fd_sc_hd__clkbuf_2 output123 (.A(net123),
    .X(eoi[29]));
 sky130_fd_sc_hd__clkbuf_2 output124 (.A(net124),
    .X(eoi[2]));
 sky130_fd_sc_hd__clkbuf_2 output125 (.A(net125),
    .X(eoi[30]));
 sky130_fd_sc_hd__clkbuf_2 output126 (.A(net126),
    .X(eoi[31]));
 sky130_fd_sc_hd__clkbuf_2 output127 (.A(net127),
    .X(eoi[3]));
 sky130_fd_sc_hd__clkbuf_2 output128 (.A(net128),
    .X(eoi[4]));
 sky130_fd_sc_hd__clkbuf_2 output129 (.A(net129),
    .X(eoi[5]));
 sky130_fd_sc_hd__clkbuf_2 output130 (.A(net130),
    .X(eoi[6]));
 sky130_fd_sc_hd__clkbuf_2 output131 (.A(net131),
    .X(eoi[7]));
 sky130_fd_sc_hd__clkbuf_2 output132 (.A(net132),
    .X(eoi[8]));
 sky130_fd_sc_hd__clkbuf_2 output133 (.A(net133),
    .X(eoi[9]));
 sky130_fd_sc_hd__clkbuf_2 output134 (.A(net134),
    .X(mem_addr[0]));
 sky130_fd_sc_hd__clkbuf_2 output135 (.A(net135),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__clkbuf_2 output136 (.A(net136),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__clkbuf_2 output137 (.A(net137),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__clkbuf_2 output138 (.A(net138),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__clkbuf_2 output139 (.A(net139),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__clkbuf_2 output140 (.A(net140),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__clkbuf_2 output141 (.A(net141),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__clkbuf_2 output142 (.A(net142),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__clkbuf_2 output143 (.A(net143),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__clkbuf_2 output144 (.A(net144),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__clkbuf_2 output145 (.A(net145),
    .X(mem_addr[1]));
 sky130_fd_sc_hd__clkbuf_2 output146 (.A(net146),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__clkbuf_2 output147 (.A(net147),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__clkbuf_2 output148 (.A(net148),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__clkbuf_2 output149 (.A(net149),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__clkbuf_2 output150 (.A(net150),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__clkbuf_2 output151 (.A(net151),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__clkbuf_2 output152 (.A(net152),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__clkbuf_2 output153 (.A(net153),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__clkbuf_2 output154 (.A(net154),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__clkbuf_2 output155 (.A(net155),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__clkbuf_2 output156 (.A(net156),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__clkbuf_2 output157 (.A(net157),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__clkbuf_2 output158 (.A(net158),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__clkbuf_2 output159 (.A(net159),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__clkbuf_2 output160 (.A(net160),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__clkbuf_2 output161 (.A(net161),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__clkbuf_2 output162 (.A(net162),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__clkbuf_2 output163 (.A(net163),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__clkbuf_2 output164 (.A(net164),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__clkbuf_2 output165 (.A(net165),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__clkbuf_2 output166 (.A(net166),
    .X(mem_instr));
 sky130_fd_sc_hd__clkbuf_2 output167 (.A(net167),
    .X(mem_la_addr[0]));
 sky130_fd_sc_hd__clkbuf_2 output168 (.A(net168),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__clkbuf_2 output169 (.A(net169),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__clkbuf_2 output170 (.A(net170),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__clkbuf_2 output171 (.A(net171),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__clkbuf_2 output172 (.A(net172),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__clkbuf_2 output173 (.A(net173),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__clkbuf_2 output174 (.A(net174),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__clkbuf_2 output175 (.A(net175),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__clkbuf_2 output176 (.A(net176),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__clkbuf_2 output177 (.A(net177),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__clkbuf_2 output178 (.A(net178),
    .X(mem_la_addr[1]));
 sky130_fd_sc_hd__clkbuf_2 output179 (.A(net179),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__clkbuf_2 output180 (.A(net180),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__clkbuf_2 output181 (.A(net181),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__clkbuf_2 output182 (.A(net182),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__clkbuf_2 output183 (.A(net183),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__clkbuf_2 output184 (.A(net184),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__clkbuf_2 output185 (.A(net185),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__clkbuf_2 output186 (.A(net186),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__clkbuf_2 output187 (.A(net187),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__clkbuf_2 output188 (.A(net188),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__clkbuf_2 output189 (.A(net189),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__clkbuf_2 output190 (.A(net190),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__clkbuf_2 output191 (.A(net191),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__clkbuf_2 output192 (.A(net192),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__clkbuf_2 output193 (.A(net193),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__clkbuf_2 output194 (.A(net194),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__clkbuf_2 output195 (.A(net195),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__clkbuf_2 output196 (.A(net196),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__clkbuf_2 output197 (.A(net197),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__clkbuf_2 output198 (.A(net198),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__clkbuf_2 output199 (.A(net199),
    .X(mem_la_read));
 sky130_fd_sc_hd__clkbuf_2 output200 (.A(net493),
    .X(mem_la_wdata[0]));
 sky130_fd_sc_hd__clkbuf_2 output201 (.A(net201),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__clkbuf_2 output202 (.A(net202),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__clkbuf_2 output203 (.A(net203),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__clkbuf_2 output204 (.A(net204),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__clkbuf_2 output205 (.A(net205),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__clkbuf_2 output206 (.A(net206),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__clkbuf_2 output207 (.A(net207),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__clkbuf_2 output208 (.A(net208),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__clkbuf_2 output209 (.A(net209),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__clkbuf_2 output210 (.A(net210),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__clkbuf_2 output211 (.A(net211),
    .X(mem_la_wdata[1]));
 sky130_fd_sc_hd__clkbuf_2 output212 (.A(net212),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__clkbuf_2 output213 (.A(net213),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__clkbuf_2 output214 (.A(net214),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__clkbuf_2 output215 (.A(net215),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__clkbuf_2 output216 (.A(net216),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__clkbuf_2 output217 (.A(net217),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__clkbuf_2 output218 (.A(net218),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__clkbuf_2 output219 (.A(net219),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__clkbuf_2 output220 (.A(net220),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__clkbuf_2 output221 (.A(net221),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__clkbuf_2 output222 (.A(net222),
    .X(mem_la_wdata[2]));
 sky130_fd_sc_hd__clkbuf_2 output223 (.A(net223),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__clkbuf_2 output224 (.A(net224),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__clkbuf_2 output225 (.A(net225),
    .X(mem_la_wdata[3]));
 sky130_fd_sc_hd__clkbuf_2 output226 (.A(net226),
    .X(mem_la_wdata[4]));
 sky130_fd_sc_hd__clkbuf_2 output227 (.A(net227),
    .X(mem_la_wdata[5]));
 sky130_fd_sc_hd__clkbuf_2 output228 (.A(net228),
    .X(mem_la_wdata[6]));
 sky130_fd_sc_hd__clkbuf_2 output229 (.A(net229),
    .X(mem_la_wdata[7]));
 sky130_fd_sc_hd__clkbuf_2 output230 (.A(net230),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__clkbuf_2 output231 (.A(net231),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__clkbuf_2 output232 (.A(net232),
    .X(mem_la_write));
 sky130_fd_sc_hd__clkbuf_2 output233 (.A(net233),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_2 output234 (.A(net234),
    .X(mem_la_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_2 output235 (.A(net235),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_2 output236 (.A(net236),
    .X(mem_la_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_2 output237 (.A(net237),
    .X(mem_valid));
 sky130_fd_sc_hd__clkbuf_2 output238 (.A(net238),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__clkbuf_2 output239 (.A(net239),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__clkbuf_2 output240 (.A(net240),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__clkbuf_2 output241 (.A(net241),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__clkbuf_2 output242 (.A(net242),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__clkbuf_2 output243 (.A(net243),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__clkbuf_2 output244 (.A(net244),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__clkbuf_2 output245 (.A(net245),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__clkbuf_2 output246 (.A(net246),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__clkbuf_2 output247 (.A(net247),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__clkbuf_2 output248 (.A(net248),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__clkbuf_2 output249 (.A(net249),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__clkbuf_2 output250 (.A(net250),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__clkbuf_2 output251 (.A(net251),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__clkbuf_2 output252 (.A(net252),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__clkbuf_2 output253 (.A(net253),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__clkbuf_2 output254 (.A(net254),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__clkbuf_2 output255 (.A(net255),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__clkbuf_2 output256 (.A(net256),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__clkbuf_2 output257 (.A(net257),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__clkbuf_2 output258 (.A(net258),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__clkbuf_2 output259 (.A(net259),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__clkbuf_2 output260 (.A(net260),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__clkbuf_2 output261 (.A(net261),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__clkbuf_2 output262 (.A(net262),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__clkbuf_2 output263 (.A(net263),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__clkbuf_2 output264 (.A(net264),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__clkbuf_2 output265 (.A(net265),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__clkbuf_2 output266 (.A(net266),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__clkbuf_2 output267 (.A(net267),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__clkbuf_2 output268 (.A(net268),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__clkbuf_2 output269 (.A(net269),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__clkbuf_2 output270 (.A(net270),
    .X(mem_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_2 output271 (.A(net271),
    .X(mem_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_2 output272 (.A(net272),
    .X(mem_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_2 output273 (.A(net273),
    .X(mem_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_2 output274 (.A(net274),
    .X(pcpi_insn[0]));
 sky130_fd_sc_hd__clkbuf_2 output275 (.A(net275),
    .X(pcpi_insn[10]));
 sky130_fd_sc_hd__clkbuf_2 output276 (.A(net276),
    .X(pcpi_insn[11]));
 sky130_fd_sc_hd__clkbuf_2 output277 (.A(net277),
    .X(pcpi_insn[12]));
 sky130_fd_sc_hd__clkbuf_2 output278 (.A(net278),
    .X(pcpi_insn[13]));
 sky130_fd_sc_hd__clkbuf_2 output279 (.A(net279),
    .X(pcpi_insn[14]));
 sky130_fd_sc_hd__clkbuf_2 output280 (.A(net280),
    .X(pcpi_insn[15]));
 sky130_fd_sc_hd__clkbuf_2 output281 (.A(net281),
    .X(pcpi_insn[16]));
 sky130_fd_sc_hd__clkbuf_2 output282 (.A(net282),
    .X(pcpi_insn[17]));
 sky130_fd_sc_hd__clkbuf_2 output283 (.A(net283),
    .X(pcpi_insn[18]));
 sky130_fd_sc_hd__clkbuf_2 output284 (.A(net284),
    .X(pcpi_insn[19]));
 sky130_fd_sc_hd__clkbuf_2 output285 (.A(net285),
    .X(pcpi_insn[1]));
 sky130_fd_sc_hd__clkbuf_2 output286 (.A(net286),
    .X(pcpi_insn[20]));
 sky130_fd_sc_hd__clkbuf_2 output287 (.A(net287),
    .X(pcpi_insn[21]));
 sky130_fd_sc_hd__clkbuf_2 output288 (.A(net288),
    .X(pcpi_insn[22]));
 sky130_fd_sc_hd__clkbuf_2 output289 (.A(net289),
    .X(pcpi_insn[23]));
 sky130_fd_sc_hd__clkbuf_2 output290 (.A(net290),
    .X(pcpi_insn[24]));
 sky130_fd_sc_hd__clkbuf_2 output291 (.A(net291),
    .X(pcpi_insn[25]));
 sky130_fd_sc_hd__clkbuf_2 output292 (.A(net292),
    .X(pcpi_insn[26]));
 sky130_fd_sc_hd__clkbuf_2 output293 (.A(net293),
    .X(pcpi_insn[27]));
 sky130_fd_sc_hd__clkbuf_2 output294 (.A(net294),
    .X(pcpi_insn[28]));
 sky130_fd_sc_hd__clkbuf_2 output295 (.A(net295),
    .X(pcpi_insn[29]));
 sky130_fd_sc_hd__clkbuf_2 output296 (.A(net296),
    .X(pcpi_insn[2]));
 sky130_fd_sc_hd__clkbuf_2 output297 (.A(net297),
    .X(pcpi_insn[30]));
 sky130_fd_sc_hd__clkbuf_2 output298 (.A(net298),
    .X(pcpi_insn[31]));
 sky130_fd_sc_hd__clkbuf_2 output299 (.A(net299),
    .X(pcpi_insn[3]));
 sky130_fd_sc_hd__clkbuf_2 output300 (.A(net300),
    .X(pcpi_insn[4]));
 sky130_fd_sc_hd__clkbuf_2 output301 (.A(net301),
    .X(pcpi_insn[5]));
 sky130_fd_sc_hd__clkbuf_2 output302 (.A(net302),
    .X(pcpi_insn[6]));
 sky130_fd_sc_hd__clkbuf_2 output303 (.A(net303),
    .X(pcpi_insn[7]));
 sky130_fd_sc_hd__clkbuf_2 output304 (.A(net304),
    .X(pcpi_insn[8]));
 sky130_fd_sc_hd__clkbuf_2 output305 (.A(net305),
    .X(pcpi_insn[9]));
 sky130_fd_sc_hd__clkbuf_2 output306 (.A(net306),
    .X(pcpi_rs1[0]));
 sky130_fd_sc_hd__clkbuf_2 output307 (.A(net307),
    .X(pcpi_rs1[10]));
 sky130_fd_sc_hd__clkbuf_2 output308 (.A(net308),
    .X(pcpi_rs1[11]));
 sky130_fd_sc_hd__clkbuf_2 output309 (.A(net309),
    .X(pcpi_rs1[12]));
 sky130_fd_sc_hd__clkbuf_2 output310 (.A(net310),
    .X(pcpi_rs1[13]));
 sky130_fd_sc_hd__clkbuf_2 output311 (.A(net311),
    .X(pcpi_rs1[14]));
 sky130_fd_sc_hd__clkbuf_2 output312 (.A(net312),
    .X(pcpi_rs1[15]));
 sky130_fd_sc_hd__clkbuf_2 output313 (.A(net313),
    .X(pcpi_rs1[16]));
 sky130_fd_sc_hd__clkbuf_2 output314 (.A(net314),
    .X(pcpi_rs1[17]));
 sky130_fd_sc_hd__clkbuf_2 output315 (.A(net315),
    .X(pcpi_rs1[18]));
 sky130_fd_sc_hd__clkbuf_2 output316 (.A(net316),
    .X(pcpi_rs1[19]));
 sky130_fd_sc_hd__clkbuf_2 output317 (.A(net317),
    .X(pcpi_rs1[1]));
 sky130_fd_sc_hd__clkbuf_2 output318 (.A(net318),
    .X(pcpi_rs1[20]));
 sky130_fd_sc_hd__clkbuf_2 output319 (.A(net319),
    .X(pcpi_rs1[21]));
 sky130_fd_sc_hd__clkbuf_2 output320 (.A(net320),
    .X(pcpi_rs1[22]));
 sky130_fd_sc_hd__clkbuf_2 output321 (.A(net321),
    .X(pcpi_rs1[23]));
 sky130_fd_sc_hd__clkbuf_2 output322 (.A(net322),
    .X(pcpi_rs1[24]));
 sky130_fd_sc_hd__clkbuf_2 output323 (.A(net323),
    .X(pcpi_rs1[25]));
 sky130_fd_sc_hd__clkbuf_2 output324 (.A(net324),
    .X(pcpi_rs1[26]));
 sky130_fd_sc_hd__clkbuf_2 output325 (.A(net325),
    .X(pcpi_rs1[27]));
 sky130_fd_sc_hd__clkbuf_2 output326 (.A(net326),
    .X(pcpi_rs1[28]));
 sky130_fd_sc_hd__clkbuf_2 output327 (.A(net327),
    .X(pcpi_rs1[29]));
 sky130_fd_sc_hd__clkbuf_2 output328 (.A(net328),
    .X(pcpi_rs1[2]));
 sky130_fd_sc_hd__clkbuf_2 output329 (.A(net329),
    .X(pcpi_rs1[30]));
 sky130_fd_sc_hd__clkbuf_2 output330 (.A(net330),
    .X(pcpi_rs1[31]));
 sky130_fd_sc_hd__clkbuf_2 output331 (.A(net331),
    .X(pcpi_rs1[3]));
 sky130_fd_sc_hd__clkbuf_2 output332 (.A(net332),
    .X(pcpi_rs1[4]));
 sky130_fd_sc_hd__clkbuf_2 output333 (.A(net333),
    .X(pcpi_rs1[5]));
 sky130_fd_sc_hd__clkbuf_2 output334 (.A(net334),
    .X(pcpi_rs1[6]));
 sky130_fd_sc_hd__clkbuf_2 output335 (.A(net335),
    .X(pcpi_rs1[7]));
 sky130_fd_sc_hd__clkbuf_2 output336 (.A(net336),
    .X(pcpi_rs1[8]));
 sky130_fd_sc_hd__clkbuf_2 output337 (.A(net337),
    .X(pcpi_rs1[9]));
 sky130_fd_sc_hd__clkbuf_2 output338 (.A(net338),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__clkbuf_2 output339 (.A(net339),
    .X(pcpi_rs2[10]));
 sky130_fd_sc_hd__clkbuf_2 output340 (.A(net340),
    .X(pcpi_rs2[11]));
 sky130_fd_sc_hd__clkbuf_2 output341 (.A(net341),
    .X(pcpi_rs2[12]));
 sky130_fd_sc_hd__clkbuf_2 output342 (.A(net342),
    .X(pcpi_rs2[13]));
 sky130_fd_sc_hd__clkbuf_2 output343 (.A(net343),
    .X(pcpi_rs2[14]));
 sky130_fd_sc_hd__clkbuf_2 output344 (.A(net344),
    .X(pcpi_rs2[15]));
 sky130_fd_sc_hd__clkbuf_2 output345 (.A(net345),
    .X(pcpi_rs2[16]));
 sky130_fd_sc_hd__clkbuf_2 output346 (.A(net346),
    .X(pcpi_rs2[17]));
 sky130_fd_sc_hd__clkbuf_2 output347 (.A(net347),
    .X(pcpi_rs2[18]));
 sky130_fd_sc_hd__clkbuf_2 output348 (.A(net348),
    .X(pcpi_rs2[19]));
 sky130_fd_sc_hd__clkbuf_2 output349 (.A(net349),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__clkbuf_2 output350 (.A(net350),
    .X(pcpi_rs2[20]));
 sky130_fd_sc_hd__clkbuf_2 output351 (.A(net351),
    .X(pcpi_rs2[21]));
 sky130_fd_sc_hd__clkbuf_2 output352 (.A(net352),
    .X(pcpi_rs2[22]));
 sky130_fd_sc_hd__clkbuf_2 output353 (.A(net353),
    .X(pcpi_rs2[23]));
 sky130_fd_sc_hd__clkbuf_2 output354 (.A(net354),
    .X(pcpi_rs2[24]));
 sky130_fd_sc_hd__clkbuf_2 output355 (.A(net355),
    .X(pcpi_rs2[25]));
 sky130_fd_sc_hd__clkbuf_2 output356 (.A(net356),
    .X(pcpi_rs2[26]));
 sky130_fd_sc_hd__clkbuf_2 output357 (.A(net357),
    .X(pcpi_rs2[27]));
 sky130_fd_sc_hd__clkbuf_2 output358 (.A(net358),
    .X(pcpi_rs2[28]));
 sky130_fd_sc_hd__clkbuf_2 output359 (.A(net359),
    .X(pcpi_rs2[29]));
 sky130_fd_sc_hd__clkbuf_2 output360 (.A(net360),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__clkbuf_2 output361 (.A(net361),
    .X(pcpi_rs2[30]));
 sky130_fd_sc_hd__clkbuf_2 output362 (.A(net362),
    .X(pcpi_rs2[31]));
 sky130_fd_sc_hd__clkbuf_2 output363 (.A(net363),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__clkbuf_2 output364 (.A(net364),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__clkbuf_2 output365 (.A(net365),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__clkbuf_2 output366 (.A(net366),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__clkbuf_2 output367 (.A(net367),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__clkbuf_2 output368 (.A(net368),
    .X(pcpi_rs2[8]));
 sky130_fd_sc_hd__clkbuf_2 output369 (.A(net369),
    .X(pcpi_rs2[9]));
 sky130_fd_sc_hd__clkbuf_2 output370 (.A(net370),
    .X(pcpi_valid));
 sky130_fd_sc_hd__clkbuf_2 output371 (.A(net371),
    .X(trace_data[0]));
 sky130_fd_sc_hd__clkbuf_2 output372 (.A(net372),
    .X(trace_data[10]));
 sky130_fd_sc_hd__clkbuf_2 output373 (.A(net373),
    .X(trace_data[11]));
 sky130_fd_sc_hd__clkbuf_2 output374 (.A(net374),
    .X(trace_data[12]));
 sky130_fd_sc_hd__clkbuf_2 output375 (.A(net375),
    .X(trace_data[13]));
 sky130_fd_sc_hd__clkbuf_2 output376 (.A(net376),
    .X(trace_data[14]));
 sky130_fd_sc_hd__clkbuf_2 output377 (.A(net377),
    .X(trace_data[15]));
 sky130_fd_sc_hd__clkbuf_2 output378 (.A(net378),
    .X(trace_data[16]));
 sky130_fd_sc_hd__clkbuf_2 output379 (.A(net379),
    .X(trace_data[17]));
 sky130_fd_sc_hd__clkbuf_2 output380 (.A(net380),
    .X(trace_data[18]));
 sky130_fd_sc_hd__clkbuf_2 output381 (.A(net381),
    .X(trace_data[19]));
 sky130_fd_sc_hd__clkbuf_2 output382 (.A(net382),
    .X(trace_data[1]));
 sky130_fd_sc_hd__clkbuf_2 output383 (.A(net383),
    .X(trace_data[20]));
 sky130_fd_sc_hd__clkbuf_2 output384 (.A(net384),
    .X(trace_data[21]));
 sky130_fd_sc_hd__clkbuf_2 output385 (.A(net385),
    .X(trace_data[22]));
 sky130_fd_sc_hd__clkbuf_2 output386 (.A(net386),
    .X(trace_data[23]));
 sky130_fd_sc_hd__clkbuf_2 output387 (.A(net387),
    .X(trace_data[24]));
 sky130_fd_sc_hd__clkbuf_2 output388 (.A(net388),
    .X(trace_data[25]));
 sky130_fd_sc_hd__clkbuf_2 output389 (.A(net389),
    .X(trace_data[26]));
 sky130_fd_sc_hd__clkbuf_2 output390 (.A(net390),
    .X(trace_data[27]));
 sky130_fd_sc_hd__clkbuf_2 output391 (.A(net391),
    .X(trace_data[28]));
 sky130_fd_sc_hd__clkbuf_2 output392 (.A(net392),
    .X(trace_data[29]));
 sky130_fd_sc_hd__clkbuf_2 output393 (.A(net393),
    .X(trace_data[2]));
 sky130_fd_sc_hd__clkbuf_2 output394 (.A(net394),
    .X(trace_data[30]));
 sky130_fd_sc_hd__clkbuf_2 output395 (.A(net395),
    .X(trace_data[31]));
 sky130_fd_sc_hd__clkbuf_2 output396 (.A(net396),
    .X(trace_data[32]));
 sky130_fd_sc_hd__clkbuf_2 output397 (.A(net397),
    .X(trace_data[33]));
 sky130_fd_sc_hd__clkbuf_2 output398 (.A(net398),
    .X(trace_data[34]));
 sky130_fd_sc_hd__clkbuf_2 output399 (.A(net399),
    .X(trace_data[35]));
 sky130_fd_sc_hd__clkbuf_2 output400 (.A(net400),
    .X(trace_data[3]));
 sky130_fd_sc_hd__clkbuf_2 output401 (.A(net401),
    .X(trace_data[4]));
 sky130_fd_sc_hd__clkbuf_2 output402 (.A(net402),
    .X(trace_data[5]));
 sky130_fd_sc_hd__clkbuf_2 output403 (.A(net403),
    .X(trace_data[6]));
 sky130_fd_sc_hd__clkbuf_2 output404 (.A(net404),
    .X(trace_data[7]));
 sky130_fd_sc_hd__clkbuf_2 output405 (.A(net405),
    .X(trace_data[8]));
 sky130_fd_sc_hd__clkbuf_2 output406 (.A(net406),
    .X(trace_data[9]));
 sky130_fd_sc_hd__clkbuf_2 output407 (.A(net407),
    .X(trace_valid));
 sky130_fd_sc_hd__clkbuf_2 output408 (.A(net408),
    .X(trap));
 sky130_fd_sc_hd__buf_4 repeater409 (.A(_09342_),
    .X(net409));
 sky130_fd_sc_hd__buf_8 repeater410 (.A(_11603_),
    .X(net410));
 sky130_fd_sc_hd__buf_8 repeater411 (.A(_12042_),
    .X(net411));
 sky130_fd_sc_hd__buf_8 repeater412 (.A(_12041_),
    .X(net412));
 sky130_fd_sc_hd__buf_6 repeater413 (.A(_10337_),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_8 repeater414 (.A(_10170_),
    .X(net414));
 sky130_fd_sc_hd__buf_6 repeater415 (.A(_11330_),
    .X(net415));
 sky130_fd_sc_hd__buf_12 repeater416 (.A(_00308_),
    .X(net416));
 sky130_fd_sc_hd__buf_4 repeater417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_6 repeater418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_4 repeater419 (.A(_01208_),
    .X(net419));
 sky130_fd_sc_hd__buf_6 repeater420 (.A(_08529_),
    .X(net420));
 sky130_fd_sc_hd__buf_12 repeater421 (.A(_02217_),
    .X(net421));
 sky130_fd_sc_hd__buf_6 repeater422 (.A(_13863_),
    .X(net422));
 sky130_fd_sc_hd__buf_6 repeater423 (.A(_13862_),
    .X(net423));
 sky130_fd_sc_hd__buf_8 repeater424 (.A(_12922_),
    .X(net424));
 sky130_fd_sc_hd__buf_6 repeater425 (.A(_12907_),
    .X(net425));
 sky130_fd_sc_hd__buf_12 repeater426 (.A(_15209_),
    .X(net426));
 sky130_fd_sc_hd__buf_8 repeater427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_8 repeater428 (.A(_14272_),
    .X(net428));
 sky130_fd_sc_hd__buf_8 repeater429 (.A(_14271_),
    .X(net429));
 sky130_fd_sc_hd__buf_8 repeater430 (.A(_14270_),
    .X(net430));
 sky130_fd_sc_hd__buf_8 repeater431 (.A(_12975_),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_8 repeater432 (.A(_12952_),
    .X(net432));
 sky130_fd_sc_hd__buf_8 repeater433 (.A(_12940_),
    .X(net433));
 sky130_fd_sc_hd__buf_8 repeater434 (.A(_12927_),
    .X(net434));
 sky130_fd_sc_hd__buf_8 repeater435 (.A(_12906_),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_8 repeater436 (.A(_01706_),
    .X(net436));
 sky130_fd_sc_hd__buf_6 repeater437 (.A(_06889_),
    .X(net437));
 sky130_fd_sc_hd__buf_6 repeater438 (.A(_05718_),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_16 repeater439 (.A(_02069_),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_8 repeater440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_8 repeater441 (.A(net443),
    .X(net441));
 sky130_fd_sc_hd__buf_6 repeater442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_8 repeater443 (.A(_00301_),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_8 repeater444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_8 repeater445 (.A(mem_xfer),
    .X(net445));
 sky130_fd_sc_hd__buf_8 repeater446 (.A(_01717_),
    .X(net446));
 sky130_fd_sc_hd__buf_8 repeater447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_8 repeater448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_12 repeater449 (.A(_00368_),
    .X(net449));
 sky130_fd_sc_hd__buf_8 repeater450 (.A(net452),
    .X(net450));
 sky130_fd_sc_hd__buf_8 repeater451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_8 repeater452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_8 repeater453 (.A(_01683_),
    .X(net453));
 sky130_fd_sc_hd__buf_8 repeater454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__buf_8 repeater455 (.A(_00292_),
    .X(net455));
 sky130_fd_sc_hd__buf_4 repeater456 (.A(_12637_),
    .X(net456));
 sky130_fd_sc_hd__buf_12 repeater457 (.A(net460),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_8 repeater458 (.A(net460),
    .X(net458));
 sky130_fd_sc_hd__buf_8 repeater459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_8 repeater460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_12 repeater461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_12 repeater462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_12 repeater463 (.A(_00357_),
    .X(net463));
 sky130_fd_sc_hd__buf_12 repeater464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_12 repeater465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_12 repeater466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_12 repeater467 (.A(_00357_),
    .X(net467));
 sky130_fd_sc_hd__buf_12 repeater468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_12 repeater469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_8 repeater470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_12 repeater471 (.A(net474),
    .X(net471));
 sky130_fd_sc_hd__buf_12 repeater472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_12 repeater473 (.A(net475),
    .X(net473));
 sky130_fd_sc_hd__buf_12 repeater474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__buf_12 repeater475 (.A(_00358_),
    .X(net475));
 sky130_fd_sc_hd__buf_12 repeater476 (.A(net478),
    .X(net476));
 sky130_fd_sc_hd__buf_12 repeater477 (.A(net478),
    .X(net477));
 sky130_fd_sc_hd__buf_12 repeater478 (.A(_00360_),
    .X(net478));
 sky130_fd_sc_hd__buf_12 repeater479 (.A(_00362_),
    .X(net479));
 sky130_fd_sc_hd__buf_12 repeater480 (.A(_00362_),
    .X(net480));
 sky130_fd_sc_hd__buf_8 repeater481 (.A(_01816_),
    .X(net481));
 sky130_fd_sc_hd__buf_8 repeater482 (.A(_01304_),
    .X(net482));
 sky130_fd_sc_hd__buf_8 repeater483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__buf_8 repeater484 (.A(_00297_),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_4 repeater485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__buf_4 repeater486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_4 repeater487 (.A(_01714_),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_16 repeater488 (.A(net226),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_16 repeater489 (.A(net225),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_16 repeater490 (.A(net222),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_16 repeater491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_16 repeater492 (.A(net211),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_16 repeater493 (.A(net200),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_16 repeater494 (.A(instr_timer),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_16 repeater495 (.A(\cpu_state[3] ),
    .X(net495));
 sky130_fd_sc_hd__buf_8 repeater496 (.A(net7),
    .X(net496));
 sky130_fd_sc_hd__buf_8 repeater497 (.A(net56),
    .X(net497));
 sky130_fd_sc_hd__buf_8 repeater498 (.A(net43),
    .X(net498));
 sky130_fd_sc_hd__buf_8 repeater499 (.A(net41),
    .X(net499));
 sky130_fd_sc_hd__buf_8 repeater500 (.A(net39),
    .X(net500));
 sky130_fd_sc_hd__buf_8 repeater501 (.A(net30),
    .X(net501));
 sky130_fd_sc_hd__buf_8 repeater502 (.A(net21),
    .X(net502));
 sky130_fd_sc_hd__buf_8 repeater503 (.A(net20),
    .X(net503));
 sky130_fd_sc_hd__buf_8 repeater504 (.A(net2),
    .X(net504));
 sky130_fd_sc_hd__buf_8 repeater505 (.A(net13),
    .X(net505));
endmodule
